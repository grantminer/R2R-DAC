magic
tech sky130A
timestamp 1700687895
<< nwell >>
rect -130 1845 3015 3120
<< nmos >>
rect -65 595 -15 1795
rect 10 595 60 1795
rect 85 595 135 1795
rect 160 595 210 1795
rect 235 595 285 1795
rect 425 595 475 1795
rect 645 595 695 1795
rect 745 595 795 1795
rect 845 595 895 1795
rect 945 595 995 1795
rect 1045 595 1095 1795
rect 1145 595 1195 1795
rect 1325 595 1375 1795
rect 1510 595 1560 1795
rect 1690 595 1740 1795
rect 1790 595 1840 1795
rect 1890 595 1940 1795
rect 1990 595 2040 1795
rect 2090 595 2140 1795
rect 2190 595 2240 1795
rect 2410 595 2460 1795
rect 2600 595 2650 1795
rect 2675 595 2725 1795
rect 2750 595 2800 1795
rect 2825 595 2875 1795
rect 2900 595 2950 1795
<< pmos >>
rect -20 1895 30 3095
rect 80 1895 130 3095
rect 180 1895 230 3095
rect 280 1895 330 3095
rect 380 1895 430 3095
rect 480 1895 530 3095
rect 660 1895 710 3095
rect 735 1895 785 3095
rect 810 1895 860 3095
rect 885 1895 935 3095
rect 960 1895 1010 3095
rect 1145 1895 1195 3095
rect 1325 1895 1375 3095
rect 1510 1895 1560 3095
rect 1690 1895 1740 3095
rect 1875 1895 1925 3095
rect 1950 1895 2000 3095
rect 2025 1895 2075 3095
rect 2100 1895 2150 3095
rect 2175 1895 2225 3095
rect 2355 1895 2405 3095
rect 2455 1895 2505 3095
rect 2555 1895 2605 3095
rect 2655 1895 2705 3095
rect 2755 1895 2805 3095
rect 2855 1895 2905 3095
<< ndiff >>
rect -115 1780 -65 1795
rect -115 610 -100 1780
rect -80 610 -65 1780
rect -115 595 -65 610
rect -15 595 10 1795
rect 60 595 85 1795
rect 135 595 160 1795
rect 210 595 235 1795
rect 285 1780 335 1795
rect 375 1780 425 1795
rect 285 610 300 1780
rect 320 610 335 1780
rect 375 610 390 1780
rect 410 610 425 1780
rect 285 595 335 610
rect 375 595 425 610
rect 475 1780 525 1795
rect 475 610 490 1780
rect 510 610 525 1780
rect 475 595 525 610
rect 600 1780 645 1795
rect 600 610 610 1780
rect 630 610 645 1780
rect 600 595 645 610
rect 695 1780 745 1795
rect 695 610 710 1780
rect 730 610 745 1780
rect 695 595 745 610
rect 795 1780 845 1795
rect 795 610 810 1780
rect 830 610 845 1780
rect 795 595 845 610
rect 895 1780 945 1795
rect 895 610 910 1780
rect 930 610 945 1780
rect 895 595 945 610
rect 995 1780 1045 1795
rect 995 610 1010 1780
rect 1030 610 1045 1780
rect 995 595 1045 610
rect 1095 1780 1145 1795
rect 1095 610 1110 1780
rect 1130 610 1145 1780
rect 1095 595 1145 610
rect 1195 1780 1245 1795
rect 1195 610 1210 1780
rect 1230 610 1245 1780
rect 1195 595 1245 610
rect 1275 1780 1325 1795
rect 1275 610 1290 1780
rect 1310 610 1325 1780
rect 1275 595 1325 610
rect 1375 1780 1420 1795
rect 1460 1780 1510 1795
rect 1375 610 1385 1780
rect 1405 610 1420 1780
rect 1460 610 1475 1780
rect 1495 610 1510 1780
rect 1375 595 1420 610
rect 1460 595 1510 610
rect 1560 1780 1610 1795
rect 1560 610 1575 1780
rect 1595 610 1610 1780
rect 1560 595 1610 610
rect 1640 1780 1690 1795
rect 1640 610 1655 1780
rect 1675 610 1690 1780
rect 1640 595 1690 610
rect 1740 1780 1790 1795
rect 1740 610 1755 1780
rect 1775 610 1790 1780
rect 1740 595 1790 610
rect 1840 1780 1890 1795
rect 1840 610 1855 1780
rect 1875 610 1890 1780
rect 1840 595 1890 610
rect 1940 1780 1990 1795
rect 1940 610 1955 1780
rect 1975 610 1990 1780
rect 1940 595 1990 610
rect 2040 1780 2090 1795
rect 2040 610 2055 1780
rect 2075 610 2090 1780
rect 2040 595 2090 610
rect 2140 1780 2190 1795
rect 2140 610 2155 1780
rect 2175 610 2190 1780
rect 2140 595 2190 610
rect 2240 1780 2285 1795
rect 2240 610 2255 1780
rect 2275 610 2285 1780
rect 2240 595 2285 610
rect 2360 1780 2410 1795
rect 2360 610 2375 1780
rect 2395 610 2410 1780
rect 2360 595 2410 610
rect 2460 1780 2510 1795
rect 2550 1780 2600 1795
rect 2460 610 2475 1780
rect 2495 610 2510 1780
rect 2550 610 2565 1780
rect 2585 610 2600 1780
rect 2460 595 2510 610
rect 2550 595 2600 610
rect 2650 595 2675 1795
rect 2725 595 2750 1795
rect 2800 595 2825 1795
rect 2875 595 2900 1795
rect 2950 1780 3000 1795
rect 2950 610 2965 1780
rect 2985 610 3000 1780
rect 2950 595 3000 610
<< pdiff >>
rect -65 3080 -20 3095
rect -65 1910 -55 3080
rect -35 1910 -20 3080
rect -65 1895 -20 1910
rect 30 3080 80 3095
rect 30 1910 45 3080
rect 65 1910 80 3080
rect 30 1895 80 1910
rect 130 3080 180 3095
rect 130 1910 145 3080
rect 165 1910 180 3080
rect 130 1895 180 1910
rect 230 3080 280 3095
rect 230 1910 245 3080
rect 265 1910 280 3080
rect 230 1895 280 1910
rect 330 3080 380 3095
rect 330 1910 345 3080
rect 365 1910 380 3080
rect 330 1895 380 1910
rect 430 3080 480 3095
rect 430 1910 445 3080
rect 465 1910 480 3080
rect 430 1895 480 1910
rect 530 3080 580 3095
rect 530 1910 545 3080
rect 565 1910 580 3080
rect 530 1895 580 1910
rect 610 3080 660 3095
rect 610 1910 625 3080
rect 645 1910 660 3080
rect 610 1895 660 1910
rect 710 1895 735 3095
rect 785 1895 810 3095
rect 860 1895 885 3095
rect 935 1895 960 3095
rect 1010 3080 1060 3095
rect 1100 3080 1145 3095
rect 1010 1910 1025 3080
rect 1045 1910 1060 3080
rect 1100 1910 1110 3080
rect 1130 1910 1145 3080
rect 1010 1895 1060 1910
rect 1100 1895 1145 1910
rect 1195 3080 1245 3095
rect 1195 1910 1210 3080
rect 1230 1910 1245 3080
rect 1195 1895 1245 1910
rect 1275 3080 1325 3095
rect 1275 1910 1290 3080
rect 1310 1910 1325 3080
rect 1275 1895 1325 1910
rect 1375 3080 1420 3095
rect 1460 3080 1510 3095
rect 1375 1910 1390 3080
rect 1410 1910 1420 3080
rect 1460 1910 1475 3080
rect 1495 1910 1510 3080
rect 1375 1895 1420 1910
rect 1460 1895 1510 1910
rect 1560 3080 1610 3095
rect 1560 1910 1575 3080
rect 1595 1910 1610 3080
rect 1560 1895 1610 1910
rect 1640 3080 1690 3095
rect 1640 1910 1655 3080
rect 1675 1910 1690 3080
rect 1640 1895 1690 1910
rect 1740 3080 1785 3095
rect 1825 3080 1875 3095
rect 1740 1910 1755 3080
rect 1775 1910 1785 3080
rect 1825 1910 1840 3080
rect 1860 1910 1875 3080
rect 1740 1895 1785 1910
rect 1825 1895 1875 1910
rect 1925 1895 1950 3095
rect 2000 1895 2025 3095
rect 2075 1895 2100 3095
rect 2150 1895 2175 3095
rect 2225 3080 2275 3095
rect 2225 1910 2240 3080
rect 2260 1910 2275 3080
rect 2225 1895 2275 1910
rect 2305 3080 2355 3095
rect 2305 1910 2320 3080
rect 2340 1910 2355 3080
rect 2305 1895 2355 1910
rect 2405 3080 2455 3095
rect 2405 1910 2420 3080
rect 2440 1910 2455 3080
rect 2405 1895 2455 1910
rect 2505 3080 2555 3095
rect 2505 1910 2520 3080
rect 2540 1910 2555 3080
rect 2505 1895 2555 1910
rect 2605 3080 2655 3095
rect 2605 1910 2620 3080
rect 2640 1910 2655 3080
rect 2605 1895 2655 1910
rect 2705 3080 2755 3095
rect 2705 1910 2720 3080
rect 2740 1910 2755 3080
rect 2705 1895 2755 1910
rect 2805 3080 2855 3095
rect 2805 1910 2820 3080
rect 2840 1910 2855 3080
rect 2805 1895 2855 1910
rect 2905 3080 2950 3095
rect 2905 1910 2920 3080
rect 2940 1910 2950 3080
rect 2905 1895 2950 1910
<< ndiffc >>
rect -100 610 -80 1780
rect 300 610 320 1780
rect 390 610 410 1780
rect 490 610 510 1780
rect 610 610 630 1780
rect 710 610 730 1780
rect 810 610 830 1780
rect 910 610 930 1780
rect 1010 610 1030 1780
rect 1110 610 1130 1780
rect 1210 610 1230 1780
rect 1290 610 1310 1780
rect 1385 610 1405 1780
rect 1475 610 1495 1780
rect 1575 610 1595 1780
rect 1655 610 1675 1780
rect 1755 610 1775 1780
rect 1855 610 1875 1780
rect 1955 610 1975 1780
rect 2055 610 2075 1780
rect 2155 610 2175 1780
rect 2255 610 2275 1780
rect 2375 610 2395 1780
rect 2475 610 2495 1780
rect 2565 610 2585 1780
rect 2965 610 2985 1780
<< pdiffc >>
rect -55 1910 -35 3080
rect 45 1910 65 3080
rect 145 1910 165 3080
rect 245 1910 265 3080
rect 345 1910 365 3080
rect 445 1910 465 3080
rect 545 1910 565 3080
rect 625 1910 645 3080
rect 1025 1910 1045 3080
rect 1110 1910 1130 3080
rect 1210 1910 1230 3080
rect 1290 1910 1310 3080
rect 1390 1910 1410 3080
rect 1475 1910 1495 3080
rect 1575 1910 1595 3080
rect 1655 1910 1675 3080
rect 1755 1910 1775 3080
rect 1840 1910 1860 3080
rect 2240 1910 2260 3080
rect 2320 1910 2340 3080
rect 2420 1910 2440 3080
rect 2520 1910 2540 3080
rect 2620 1910 2640 3080
rect 2720 1910 2740 3080
rect 2820 1910 2840 3080
rect 2920 1910 2940 3080
<< psubdiff >>
rect 335 1780 375 1795
rect 335 610 345 1780
rect 365 610 375 1780
rect 335 595 375 610
rect 555 1780 600 1795
rect 555 610 570 1780
rect 590 610 600 1780
rect 555 595 600 610
rect 1420 1780 1460 1795
rect 1420 610 1430 1780
rect 1450 610 1460 1780
rect 1420 595 1460 610
rect 2285 1780 2330 1795
rect 2285 610 2295 1780
rect 2315 610 2330 1780
rect 2285 595 2330 610
rect 2510 1780 2550 1795
rect 2510 610 2520 1780
rect 2540 610 2550 1780
rect 2510 595 2550 610
<< nsubdiff >>
rect -110 3080 -65 3095
rect -110 1910 -95 3080
rect -75 1910 -65 3080
rect -110 1895 -65 1910
rect 1060 3080 1100 3095
rect 1060 1910 1070 3080
rect 1090 1910 1100 3080
rect 1060 1895 1100 1910
rect 1420 3080 1460 3095
rect 1420 1910 1430 3080
rect 1450 1910 1460 3080
rect 1420 1895 1460 1910
rect 1785 3080 1825 3095
rect 1785 1910 1795 3080
rect 1815 1910 1825 3080
rect 1785 1895 1825 1910
rect 2950 3080 2995 3095
rect 2950 1910 2960 3080
rect 2980 1910 2995 3080
rect 2950 1895 2995 1910
<< psubdiffcont >>
rect 345 610 365 1780
rect 570 610 590 1780
rect 1430 610 1450 1780
rect 2295 610 2315 1780
rect 2520 610 2540 1780
<< nsubdiffcont >>
rect -95 1910 -75 3080
rect 1070 1910 1090 3080
rect 1430 1910 1450 3080
rect 1795 1910 1815 3080
rect 2960 1910 2980 3080
<< poly >>
rect 1145 3255 1195 3260
rect 1145 3235 1160 3255
rect 1180 3235 1195 3255
rect 1145 3150 1195 3235
rect 660 3135 1195 3150
rect -20 3095 30 3110
rect 80 3095 130 3110
rect 180 3095 230 3110
rect 280 3095 330 3110
rect 380 3095 430 3110
rect 480 3095 530 3110
rect 660 3095 710 3135
rect 735 3095 785 3135
rect 810 3095 860 3135
rect 885 3095 935 3135
rect 960 3095 1010 3135
rect 1145 3095 1195 3135
rect 1325 3255 1375 3260
rect 1325 3235 1340 3255
rect 1360 3235 1375 3255
rect 1325 3095 1375 3235
rect 1510 3255 1560 3260
rect 1510 3235 1525 3255
rect 1545 3235 1560 3255
rect 1510 3095 1560 3235
rect 1690 3255 1740 3260
rect 1690 3235 1705 3255
rect 1725 3235 1740 3255
rect 1690 3150 1740 3235
rect 1690 3135 2225 3150
rect 1690 3095 1740 3135
rect 1875 3095 1925 3135
rect 1950 3095 2000 3135
rect 2025 3095 2075 3135
rect 2100 3095 2150 3135
rect 2175 3095 2225 3135
rect 2355 3095 2405 3110
rect 2455 3095 2505 3110
rect 2555 3095 2605 3110
rect 2655 3095 2705 3110
rect 2755 3095 2805 3110
rect 2855 3095 2905 3110
rect -115 1870 -65 1875
rect -115 1850 -100 1870
rect -80 1860 -65 1870
rect -20 1860 30 1895
rect 80 1875 130 1895
rect 180 1875 230 1895
rect 80 1870 230 1875
rect 80 1860 145 1870
rect -80 1850 145 1860
rect 165 1860 230 1870
rect 280 1875 330 1895
rect 380 1875 430 1895
rect 280 1870 430 1875
rect 280 1860 345 1870
rect 165 1850 345 1860
rect 365 1850 430 1870
rect -115 1845 430 1850
rect 480 1875 530 1895
rect 660 1880 710 1895
rect 735 1880 785 1895
rect 810 1880 860 1895
rect 885 1880 935 1895
rect 960 1880 1010 1895
rect 1145 1880 1195 1895
rect 1325 1880 1375 1895
rect 1510 1880 1560 1895
rect 1690 1880 1740 1895
rect 1875 1880 1925 1895
rect 1950 1880 2000 1895
rect 2025 1880 2075 1895
rect 2100 1880 2150 1895
rect 2175 1880 2225 1895
rect 2355 1875 2405 1895
rect 480 1870 580 1875
rect 480 1850 545 1870
rect 565 1850 580 1870
rect 2305 1870 2405 1875
rect 480 1845 580 1850
rect 610 1850 695 1855
rect 610 1830 625 1850
rect 645 1830 695 1850
rect 610 1825 695 1830
rect -65 1795 -15 1810
rect 10 1795 60 1810
rect 85 1795 135 1810
rect 160 1795 210 1810
rect 235 1795 285 1810
rect 425 1795 475 1810
rect 645 1795 695 1825
rect 2190 1850 2275 1855
rect 2190 1830 2240 1850
rect 2260 1830 2275 1850
rect 2305 1850 2320 1870
rect 2340 1850 2405 1870
rect 2305 1845 2405 1850
rect 2455 1875 2505 1895
rect 2555 1875 2605 1895
rect 2455 1870 2605 1875
rect 2455 1850 2520 1870
rect 2540 1860 2605 1870
rect 2655 1875 2705 1895
rect 2755 1875 2805 1895
rect 2655 1870 2805 1875
rect 2655 1860 2720 1870
rect 2540 1850 2720 1860
rect 2740 1860 2805 1870
rect 2855 1860 2905 1895
rect 2950 1870 3000 1875
rect 2950 1860 2965 1870
rect 2740 1850 2965 1860
rect 2985 1850 3000 1870
rect 2455 1845 3000 1850
rect 2190 1825 2275 1830
rect 745 1795 795 1810
rect 845 1795 895 1810
rect 945 1795 995 1810
rect 1045 1795 1095 1810
rect 1145 1795 1195 1810
rect 1325 1795 1375 1810
rect 1510 1795 1560 1810
rect 1690 1795 1740 1810
rect 1790 1795 1840 1810
rect 1890 1795 1940 1810
rect 1990 1795 2040 1810
rect 2090 1795 2140 1810
rect 2190 1795 2240 1825
rect 2410 1795 2460 1810
rect 2600 1795 2650 1810
rect 2675 1795 2725 1810
rect 2750 1795 2800 1810
rect 2825 1795 2875 1810
rect 2900 1795 2950 1810
rect -65 565 -15 595
rect 10 565 60 595
rect 85 565 135 595
rect 160 565 210 595
rect 235 565 285 595
rect 425 565 475 595
rect -65 550 475 565
rect 425 470 475 550
rect 645 560 695 595
rect 745 575 795 595
rect 845 575 895 595
rect 745 570 895 575
rect 745 560 810 570
rect 645 550 810 560
rect 830 560 895 570
rect 945 575 995 595
rect 1045 575 1095 595
rect 945 570 1095 575
rect 945 560 1010 570
rect 830 550 1010 560
rect 1030 550 1095 570
rect 645 545 1095 550
rect 1145 580 1195 595
rect 1145 575 1245 580
rect 1145 555 1210 575
rect 1230 555 1245 575
rect 1145 550 1245 555
rect 1325 575 1375 595
rect 1325 555 1340 575
rect 1360 555 1375 575
rect 1325 550 1375 555
rect 1510 575 1560 595
rect 1690 580 1740 595
rect 1510 555 1525 575
rect 1545 555 1560 575
rect 1510 550 1560 555
rect 1640 575 1740 580
rect 1640 555 1655 575
rect 1675 555 1740 575
rect 1640 550 1740 555
rect 1145 525 1195 550
rect 1690 525 1740 550
rect 1790 575 1840 595
rect 1890 575 1940 595
rect 1790 570 1940 575
rect 1790 550 1855 570
rect 1875 560 1940 570
rect 1990 575 2040 595
rect 2090 575 2140 595
rect 1990 570 2140 575
rect 1990 560 2055 570
rect 1875 550 2055 560
rect 2075 560 2140 570
rect 2190 560 2240 595
rect 2075 550 2240 560
rect 1790 545 2240 550
rect 2410 565 2460 595
rect 2600 565 2650 595
rect 2675 565 2725 595
rect 2750 565 2800 595
rect 2825 565 2875 595
rect 2900 565 2950 595
rect 2410 550 2950 565
rect 1145 500 1740 525
rect 425 450 440 470
rect 460 450 475 470
rect 425 445 475 450
rect 2410 470 2460 550
rect 2410 450 2425 470
rect 2445 450 2460 470
rect 2410 445 2460 450
<< polycont >>
rect 1160 3235 1180 3255
rect 1340 3235 1360 3255
rect 1525 3235 1545 3255
rect 1705 3235 1725 3255
rect -100 1850 -80 1870
rect 145 1850 165 1870
rect 345 1850 365 1870
rect 545 1850 565 1870
rect 625 1830 645 1850
rect 2240 1830 2260 1850
rect 2320 1850 2340 1870
rect 2520 1850 2540 1870
rect 2720 1850 2740 1870
rect 2965 1850 2985 1870
rect 810 550 830 570
rect 1010 550 1030 570
rect 1210 555 1230 575
rect 1340 555 1360 575
rect 1525 555 1545 575
rect 1655 555 1675 575
rect 1855 550 1875 570
rect 2055 550 2075 570
rect 440 450 460 470
rect 2425 450 2445 470
<< locali >>
rect -225 3255 1740 3260
rect -225 3235 1160 3255
rect 1180 3235 1340 3255
rect 1360 3235 1525 3255
rect 1545 3235 1705 3255
rect 1725 3235 1740 3255
rect -225 3230 1740 3235
rect 535 3170 3090 3200
rect 35 3110 480 3145
rect -105 3090 -65 3100
rect -105 3080 -25 3090
rect -105 1910 -95 3080
rect -75 1910 -55 3080
rect -35 1910 -25 3080
rect -105 1900 -25 1910
rect 35 3080 75 3110
rect 35 1910 45 3080
rect 65 1910 75 3080
rect 35 1900 75 1910
rect 135 3080 175 3090
rect 135 1910 145 3080
rect 165 1910 175 3080
rect 135 1875 175 1910
rect 235 3080 275 3110
rect 235 1910 245 3080
rect 265 1910 275 3080
rect 235 1900 275 1910
rect 335 3080 375 3090
rect 335 1910 345 3080
rect 365 1910 375 3080
rect 335 1875 375 1910
rect 435 3080 480 3110
rect 435 1910 445 3080
rect 465 1910 480 3080
rect 435 1900 480 1910
rect 535 3080 575 3170
rect 535 1910 545 3080
rect 565 1910 575 3080
rect 535 1875 575 1910
rect 615 3080 655 3090
rect 615 1910 625 3080
rect 645 1910 655 3080
rect -115 1870 -65 1875
rect -115 1850 -100 1870
rect -80 1850 -65 1870
rect -115 1845 -65 1850
rect 130 1870 180 1875
rect 130 1850 145 1870
rect 165 1850 180 1870
rect 130 1845 180 1850
rect 330 1870 380 1875
rect 330 1850 345 1870
rect 365 1850 380 1870
rect 330 1845 380 1850
rect 480 1870 580 1875
rect 480 1850 545 1870
rect 565 1850 580 1870
rect 615 1855 655 1910
rect 1015 3080 1140 3090
rect 1015 1910 1025 3080
rect 1045 1910 1070 3080
rect 1090 1910 1110 3080
rect 1130 1910 1140 3080
rect 1015 1900 1140 1910
rect 1200 3080 1240 3090
rect 1200 1910 1210 3080
rect 1230 1910 1240 3080
rect 480 1845 580 1850
rect 610 1850 660 1855
rect -110 1780 -70 1845
rect -110 610 -100 1780
rect -80 610 -70 1780
rect -110 600 -70 610
rect 290 1780 420 1790
rect 290 610 300 1780
rect 325 610 345 1780
rect 365 610 385 1780
rect 410 610 420 1780
rect 290 600 420 610
rect 480 1780 520 1845
rect 610 1830 625 1850
rect 645 1830 660 1850
rect 610 1825 660 1830
rect 700 1810 1145 1845
rect 480 610 490 1780
rect 510 610 520 1780
rect 480 600 520 610
rect 560 1780 640 1790
rect 560 610 570 1780
rect 590 610 610 1780
rect 630 610 640 1780
rect 560 600 640 610
rect 700 1780 740 1810
rect 700 610 710 1780
rect 730 610 740 1780
rect 700 600 740 610
rect 800 1780 840 1790
rect 800 610 810 1780
rect 830 610 840 1780
rect 800 575 840 610
rect 900 1780 940 1810
rect 900 610 910 1780
rect 930 610 940 1780
rect 900 600 940 610
rect 1000 1780 1040 1790
rect 1000 610 1010 1780
rect 1030 610 1040 1780
rect 1000 575 1040 610
rect 1100 1780 1145 1810
rect 1100 610 1110 1780
rect 1130 610 1145 1780
rect 1100 600 1145 610
rect 1200 1780 1240 1910
rect 1200 610 1210 1780
rect 1230 610 1240 1780
rect 1200 580 1240 610
rect 1280 3080 1320 3090
rect 1280 1910 1290 3080
rect 1310 1910 1320 3080
rect 1280 1780 1320 1910
rect 1375 3080 1505 3090
rect 1375 1910 1390 3080
rect 1410 1910 1430 3080
rect 1450 1910 1475 3080
rect 1495 1910 1505 3080
rect 1375 1900 1505 1910
rect 1565 3080 1605 3090
rect 1565 1910 1575 3080
rect 1595 1910 1605 3080
rect 1280 610 1290 1780
rect 1310 610 1320 1780
rect 1280 580 1320 610
rect 1375 1780 1505 1790
rect 1375 610 1385 1780
rect 1410 610 1430 1780
rect 1450 610 1470 1780
rect 1495 610 1505 1780
rect 1375 600 1505 610
rect 1565 1780 1605 1910
rect 1565 610 1575 1780
rect 1595 610 1605 1780
rect 1565 580 1605 610
rect 1645 3080 1685 3090
rect 1645 1910 1655 3080
rect 1675 1910 1685 3080
rect 1645 1780 1685 1910
rect 1745 3080 1870 3090
rect 1745 1910 1755 3080
rect 1775 1910 1795 3080
rect 1815 1910 1840 3080
rect 1860 1910 1870 3080
rect 1745 1900 1870 1910
rect 2230 3080 2270 3090
rect 2230 1910 2240 3080
rect 2260 1910 2270 3080
rect 2230 1855 2270 1910
rect 2310 3080 2350 3170
rect 2310 1910 2320 3080
rect 2340 1910 2350 3080
rect 2310 1875 2350 1910
rect 2405 3110 2850 3145
rect 2405 3080 2450 3110
rect 2405 1910 2420 3080
rect 2440 1910 2450 3080
rect 2405 1900 2450 1910
rect 2510 3080 2550 3090
rect 2510 1910 2520 3080
rect 2540 1910 2550 3080
rect 2510 1875 2550 1910
rect 2610 3080 2650 3110
rect 2610 1910 2620 3080
rect 2640 1910 2650 3080
rect 2610 1900 2650 1910
rect 2710 3080 2750 3090
rect 2710 1910 2720 3080
rect 2740 1910 2750 3080
rect 2710 1875 2750 1910
rect 2810 3080 2850 3110
rect 2950 3090 2990 3100
rect 2810 1910 2820 3080
rect 2840 1910 2850 3080
rect 2810 1900 2850 1910
rect 2910 3080 2990 3090
rect 2910 1910 2920 3080
rect 2940 1910 2960 3080
rect 2980 1910 2990 3080
rect 2910 1900 2990 1910
rect 2305 1870 2405 1875
rect 2225 1850 2275 1855
rect 1645 610 1655 1780
rect 1675 610 1685 1780
rect 1645 580 1685 610
rect 1740 1810 2185 1845
rect 2225 1830 2240 1850
rect 2260 1830 2275 1850
rect 2305 1850 2320 1870
rect 2340 1850 2405 1870
rect 2305 1845 2405 1850
rect 2505 1870 2555 1875
rect 2505 1850 2520 1870
rect 2540 1850 2555 1870
rect 2505 1845 2555 1850
rect 2705 1870 2755 1875
rect 2705 1850 2720 1870
rect 2740 1850 2755 1870
rect 2705 1845 2755 1850
rect 2950 1870 3000 1875
rect 2950 1850 2965 1870
rect 2985 1850 3000 1870
rect 2950 1845 3000 1850
rect 2225 1825 2275 1830
rect 1740 1780 1785 1810
rect 1740 610 1755 1780
rect 1775 610 1785 1780
rect 1740 600 1785 610
rect 1845 1780 1885 1790
rect 1845 610 1855 1780
rect 1875 610 1885 1780
rect 1195 575 1245 580
rect 795 570 845 575
rect 795 550 810 570
rect 830 550 845 570
rect 795 545 845 550
rect 995 570 1045 575
rect 995 550 1010 570
rect 1030 550 1045 570
rect 1195 555 1210 575
rect 1230 555 1245 575
rect 1195 550 1245 555
rect 1280 575 1375 580
rect 1280 555 1340 575
rect 1360 555 1375 575
rect 1280 550 1375 555
rect 995 545 1045 550
rect 425 470 475 475
rect 1325 470 1375 550
rect 1510 575 1605 580
rect 1510 555 1525 575
rect 1545 555 1605 575
rect 1510 550 1605 555
rect 1640 575 1690 580
rect 1845 575 1885 610
rect 1945 1780 1985 1810
rect 1945 610 1955 1780
rect 1975 610 1985 1780
rect 1945 600 1985 610
rect 2045 1780 2085 1790
rect 2045 610 2055 1780
rect 2075 610 2085 1780
rect 2045 575 2085 610
rect 2145 1780 2185 1810
rect 2145 610 2155 1780
rect 2175 610 2185 1780
rect 2145 600 2185 610
rect 2245 1780 2325 1790
rect 2245 610 2255 1780
rect 2275 610 2295 1780
rect 2315 610 2325 1780
rect 2245 600 2325 610
rect 2365 1780 2405 1845
rect 2365 610 2375 1780
rect 2395 610 2405 1780
rect 2365 600 2405 610
rect 2465 1780 2595 1790
rect 2465 610 2475 1780
rect 2500 610 2520 1780
rect 2540 610 2560 1780
rect 2585 610 2595 1780
rect 2465 600 2595 610
rect 2955 1780 2995 1845
rect 2955 610 2965 1780
rect 2985 610 2995 1780
rect 2955 600 2995 610
rect 3016 1220 3085 1250
rect 1640 555 1655 575
rect 1675 555 1690 575
rect 1510 470 1560 550
rect 1640 520 1690 555
rect 1840 570 1890 575
rect 1840 550 1855 570
rect 1875 550 1890 570
rect 1840 545 1890 550
rect 2040 570 2090 575
rect 2040 550 2055 570
rect 2075 550 2090 570
rect 2040 545 2090 550
rect 3016 520 3041 1220
rect 1640 495 3041 520
rect 2410 470 2460 475
rect 425 450 440 470
rect 460 450 2425 470
rect 2445 450 2460 470
rect 425 445 2460 450
<< viali >>
rect -95 1910 -75 3080
rect -55 1910 -35 3080
rect 1025 1910 1045 3080
rect 1070 1910 1090 3080
rect 1110 1910 1130 3080
rect 300 610 320 1780
rect 320 610 325 1780
rect 345 610 365 1780
rect 385 610 390 1780
rect 390 610 410 1780
rect 570 610 590 1780
rect 610 610 630 1780
rect 1390 1910 1410 3080
rect 1430 1910 1450 3080
rect 1475 1910 1495 3080
rect 1385 610 1405 1780
rect 1405 610 1410 1780
rect 1430 610 1450 1780
rect 1470 610 1475 1780
rect 1475 610 1495 1780
rect 1755 1910 1775 3080
rect 1795 1910 1815 3080
rect 1840 1910 1860 3080
rect 2920 1910 2940 3080
rect 2960 1910 2980 3080
rect 2255 610 2275 1780
rect 2295 610 2315 1780
rect 2475 610 2495 1780
rect 2495 610 2500 1780
rect 2520 610 2540 1780
rect 2560 610 2565 1780
rect 2565 610 2585 1780
<< metal1 >>
rect -200 3080 3085 3095
rect -200 1910 -95 3080
rect -75 1910 -55 3080
rect -35 1910 1025 3080
rect 1045 1910 1070 3080
rect 1090 1910 1110 3080
rect 1130 1910 1390 3080
rect 1410 1910 1430 3080
rect 1450 1910 1475 3080
rect 1495 1910 1755 3080
rect 1775 1910 1795 3080
rect 1815 1910 1840 3080
rect 1860 1910 2920 3080
rect 2940 1910 2960 3080
rect 2980 1910 3085 3080
rect -200 1895 3085 1910
rect -200 1780 3085 1795
rect -200 610 300 1780
rect 325 610 345 1780
rect 365 610 385 1780
rect 410 610 570 1780
rect 590 610 610 1780
rect 630 610 1385 1780
rect 1410 610 1430 1780
rect 1450 610 1470 1780
rect 1495 610 2255 1780
rect 2275 610 2295 1780
rect 2315 610 2475 1780
rect 2500 610 2520 1780
rect 2540 610 2560 1780
rect 2585 610 3085 1780
rect -200 595 3085 610
<< labels >>
rlabel metal1 -200 2725 -200 2725 7 VP
port 3 w
rlabel locali 3085 1235 3085 1235 3 Vcn
port 5 w
rlabel metal1 -200 1185 -200 1185 7 VN
port 9 w
rlabel locali 3090 3185 3090 3185 3 Vcp
port 2 w
rlabel locali -225 3245 -225 3245 7 Vbp
port 1 w
<< end >>
