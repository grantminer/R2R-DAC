magic
tech sky130A
timestamp 1701110497
<< nwell >>
rect 1000 4905 1435 4925
rect 160 4900 4130 4905
rect 160 4899 5650 4900
rect 160 3660 5705 4899
rect 220 2990 5705 3660
rect 160 1750 5705 2990
rect 160 1745 3890 1750
rect 5506 1749 5705 1750
rect 940 1720 1450 1745
<< nmos >>
rect 450 5145 850 6345
rect 2040 5145 2440 6345
rect 3270 5145 3670 6345
rect 4860 5145 5260 6345
rect 450 385 850 1585
rect 2040 385 2440 1585
rect 3270 385 3670 1585
rect 4860 385 5260 1585
<< pmos >>
rect 580 3680 980 4880
rect 1380 3680 1780 4880
rect 2610 3680 3010 4880
rect 3410 3680 3805 4880
rect 4645 3680 5045 4880
rect 580 1770 980 2970
rect 1380 1770 1780 2970
rect 2610 1770 3010 2970
rect 3410 1770 3805 2970
rect 4645 1770 5045 2970
<< ndiff >>
rect 50 6285 450 6345
rect 50 5205 110 6285
rect 390 5205 450 6285
rect 50 5145 450 5205
rect 850 6285 1250 6345
rect 1640 6285 2040 6345
rect 850 5205 910 6285
rect 1190 5205 1250 6285
rect 1640 5205 1700 6285
rect 1980 5205 2040 6285
rect 850 5145 1250 5205
rect 1640 5145 2040 5205
rect 2440 6285 2840 6345
rect 2440 5205 2500 6285
rect 2780 5205 2840 6285
rect 2440 5145 2840 5205
rect 2870 6285 3270 6345
rect 2870 5205 2930 6285
rect 3210 5205 3270 6285
rect 2870 5145 3270 5205
rect 3670 6285 4070 6345
rect 4460 6285 4860 6345
rect 3670 5205 3730 6285
rect 4010 5205 4070 6285
rect 4460 5205 4520 6285
rect 4800 5205 4860 6285
rect 3670 5145 4070 5205
rect 4460 5145 4860 5205
rect 5260 6285 5660 6345
rect 5260 5205 5320 6285
rect 5600 5205 5660 6285
rect 5260 5145 5660 5205
rect 50 1525 450 1585
rect 50 445 110 1525
rect 390 445 450 1525
rect 50 385 450 445
rect 850 1525 1250 1585
rect 1640 1525 2040 1585
rect 850 445 910 1525
rect 1190 445 1250 1525
rect 1640 445 1700 1525
rect 1980 445 2040 1525
rect 850 385 1250 445
rect 1640 385 2040 445
rect 2440 1525 2840 1585
rect 2440 445 2500 1525
rect 2780 445 2840 1525
rect 2440 385 2840 445
rect 2870 1525 3270 1585
rect 2870 445 2930 1525
rect 3210 445 3270 1525
rect 2870 385 3270 445
rect 3670 1525 4070 1585
rect 4460 1525 4860 1585
rect 3670 445 3730 1525
rect 4010 445 4070 1525
rect 4460 445 4520 1525
rect 4800 445 4860 1525
rect 3670 385 4070 445
rect 4460 385 4860 445
rect 5260 1525 5660 1585
rect 5260 445 5320 1525
rect 5600 445 5660 1525
rect 5260 385 5660 445
<< pdiff >>
rect 180 4820 580 4880
rect 180 3740 240 4820
rect 520 3740 580 4820
rect 180 3680 580 3740
rect 980 4820 1380 4880
rect 980 3740 1040 4820
rect 1320 3740 1380 4820
rect 980 3680 1380 3740
rect 1780 4820 2180 4880
rect 1780 3740 1840 4820
rect 2120 3740 2180 4820
rect 1780 3680 2180 3740
rect 2210 4820 2610 4880
rect 2210 3740 2270 4820
rect 2550 3740 2610 4820
rect 2210 3680 2610 3740
rect 3010 4820 3410 4880
rect 3010 3740 3070 4820
rect 3350 3740 3410 4820
rect 3010 3680 3410 3740
rect 3805 4820 4205 4880
rect 3805 3740 3865 4820
rect 4145 3740 4205 4820
rect 3805 3680 4205 3740
rect 4245 4820 4645 4880
rect 4245 3740 4305 4820
rect 4585 3740 4645 4820
rect 4245 3680 4645 3740
rect 5045 4820 5445 4880
rect 5045 3740 5105 4820
rect 5385 3740 5445 4820
rect 5045 3680 5445 3740
rect 180 2910 580 2970
rect 180 1830 240 2910
rect 520 1830 580 2910
rect 180 1770 580 1830
rect 980 2910 1380 2970
rect 980 1830 1040 2910
rect 1320 1830 1380 2910
rect 980 1770 1380 1830
rect 1780 2910 2180 2970
rect 1780 1830 1840 2910
rect 2120 1830 2180 2910
rect 1780 1770 2180 1830
rect 2210 2910 2610 2970
rect 2210 1830 2270 2910
rect 2550 1830 2610 2910
rect 2210 1770 2610 1830
rect 3010 2910 3410 2970
rect 3010 1830 3070 2910
rect 3350 1830 3410 2910
rect 3010 1770 3410 1830
rect 3805 2910 4205 2970
rect 3805 1830 3865 2910
rect 4145 1830 4205 2910
rect 3805 1770 4205 1830
rect 4245 2910 4645 2970
rect 4245 1830 4305 2910
rect 4585 1830 4645 2910
rect 4245 1770 4645 1830
rect 5045 2910 5445 2970
rect 5045 1830 5105 2910
rect 5385 1830 5445 2910
rect 5045 1770 5445 1830
<< ndiffc >>
rect 110 5205 390 6285
rect 910 5205 1190 6285
rect 1700 5205 1980 6285
rect 2500 5205 2780 6285
rect 2930 5205 3210 6285
rect 3730 5205 4010 6285
rect 4520 5205 4800 6285
rect 5320 5205 5600 6285
rect 110 445 390 1525
rect 910 445 1190 1525
rect 1700 445 1980 1525
rect 2500 445 2780 1525
rect 2930 445 3210 1525
rect 3730 445 4010 1525
rect 4520 445 4800 1525
rect 5320 445 5600 1525
<< pdiffc >>
rect 240 3740 520 4820
rect 1040 3740 1320 4820
rect 1840 3740 2120 4820
rect 2270 3740 2550 4820
rect 3070 3740 3350 4820
rect 3865 3740 4145 4820
rect 4305 3740 4585 4820
rect 5105 3740 5385 4820
rect 240 1830 520 2910
rect 1040 1830 1320 2910
rect 1840 1830 2120 2910
rect 2270 1830 2550 2910
rect 3070 1830 3350 2910
rect 3865 1830 4145 2910
rect 4305 1830 4585 2910
rect 5105 1830 5385 2910
<< psubdiff >>
rect 1250 6285 1640 6345
rect 1250 5205 1305 6285
rect 1585 5205 1640 6285
rect 1250 5145 1640 5205
rect 4070 6285 4460 6345
rect 4070 5205 4125 6285
rect 4405 5205 4460 6285
rect 4070 5145 4460 5205
rect 1250 1525 1640 1585
rect 1250 445 1305 1525
rect 1585 445 1640 1525
rect 1250 385 1640 445
rect 4070 1525 4460 1585
rect 4070 445 4125 1525
rect 4405 445 4460 1525
rect 4070 385 4460 445
<< nsubdiff >>
rect 715 3465 1915 3520
rect 715 3185 775 3465
rect 1855 3185 1915 3465
rect 715 3130 1915 3185
rect 2550 3465 3750 3520
rect 2550 3185 2610 3465
rect 3690 3185 3750 3465
rect 2550 3135 3750 3185
rect 4050 3465 5250 3520
rect 4050 3185 4110 3465
rect 5190 3185 5250 3465
rect 4050 3135 5250 3185
<< psubdiffcont >>
rect 1305 5205 1585 6285
rect 4125 5205 4405 6285
rect 1305 445 1585 1525
rect 4125 445 4405 1525
<< nsubdiffcont >>
rect 775 3185 1855 3465
rect 2610 3185 3690 3465
rect 4110 3185 5190 3465
<< poly >>
rect 450 6345 850 6375
rect 2040 6345 2440 6375
rect 3270 6345 3670 6375
rect 4860 6345 5260 6375
rect 450 5135 850 5145
rect 450 5125 1070 5135
rect 450 5105 1040 5125
rect 1060 5115 1070 5125
rect 2040 5115 2440 5145
rect 1060 5105 2440 5115
rect 450 5095 2440 5105
rect 3270 5115 3670 5145
rect 4860 5135 5260 5145
rect 4860 5125 5480 5135
rect 4860 5115 5450 5125
rect 3270 5105 5450 5115
rect 5470 5105 5480 5125
rect 3270 5100 5480 5105
rect 5440 5095 5480 5100
rect 1955 4960 1995 4970
rect 1380 4940 1965 4960
rect 1985 4940 3010 4960
rect 1380 4930 3010 4940
rect 580 4880 980 4930
rect 1380 4880 1780 4930
rect 2610 4880 3010 4930
rect 3410 4880 3805 4930
rect 4645 4880 5045 4930
rect 580 3590 980 3680
rect 1380 3630 1780 3680
rect 2610 3630 3010 3680
rect 3410 3590 3805 3680
rect 4645 3590 5045 3680
rect 580 3585 5045 3590
rect 580 3580 5475 3585
rect 580 3560 2395 3580
rect 2415 3560 5475 3580
rect 580 3540 5475 3560
rect 5400 3145 5475 3540
rect 5643 3145 5705 3146
rect 5400 3110 5705 3145
rect 580 3090 5705 3110
rect 580 3070 2395 3090
rect 2415 3087 5705 3090
rect 2415 3070 5675 3087
rect 580 3065 5675 3070
rect 580 3060 5045 3065
rect 580 2970 980 3060
rect 3405 3055 3805 3060
rect 1380 2970 1780 3020
rect 2610 2970 3010 3020
rect 3410 2970 3805 3055
rect 4645 2970 5045 3060
rect 5665 3027 5675 3065
rect 5695 3027 5705 3087
rect 5665 3017 5705 3027
rect 580 1720 980 1770
rect 1380 1720 1780 1770
rect 2610 1720 3010 1770
rect 3410 1720 3805 1770
rect 4645 1720 5045 1770
rect 1380 1710 3010 1720
rect 1380 1690 1965 1710
rect 1985 1690 3010 1710
rect 1955 1680 1995 1690
rect 450 1625 2440 1635
rect 5440 1630 5480 1635
rect 450 1605 1040 1625
rect 1060 1615 2440 1625
rect 1060 1605 1070 1615
rect 450 1595 1070 1605
rect 450 1585 850 1595
rect 2040 1585 2440 1615
rect 3270 1625 5480 1630
rect 3270 1615 5450 1625
rect 3270 1585 3670 1615
rect 4860 1605 5450 1615
rect 5470 1605 5480 1625
rect 4860 1595 5480 1605
rect 4860 1585 5260 1595
rect 450 355 850 385
rect 2040 355 2440 385
rect 3270 355 3670 385
rect 4860 355 5260 385
<< polycont >>
rect 1040 5105 1060 5125
rect 5450 5105 5470 5125
rect 1965 4940 1985 4960
rect 2395 3560 2415 3580
rect 2395 3070 2415 3090
rect 5675 3027 5695 3087
rect 1965 1690 1985 1710
rect 1040 1605 1060 1625
rect 5450 1605 5470 1625
<< locali >>
rect 80 6285 420 6320
rect 80 5205 110 6285
rect 390 5205 420 6285
rect 80 5175 420 5205
rect 880 6285 1220 6315
rect 880 5205 910 6285
rect 1190 5205 1220 6285
rect 880 5175 1220 5205
rect 1275 6285 2010 6315
rect 1275 5205 1300 6285
rect 1585 5205 1695 6285
rect 1980 5205 2010 6285
rect 1275 5175 2010 5205
rect 2470 6285 2810 6315
rect 2470 5205 2500 6285
rect 2780 5205 2810 6285
rect 2470 5175 2810 5205
rect 2900 6285 3240 6315
rect 2900 5205 2930 6285
rect 3210 5205 3240 6285
rect 2900 5175 3240 5205
rect 3700 6285 4830 6315
rect 3700 5205 3730 6285
rect 4015 5205 4120 6285
rect 4405 5205 4520 6285
rect 4805 5205 4830 6285
rect 3700 5175 4830 5205
rect 5290 6285 5630 6315
rect 5290 5205 5320 6285
rect 5600 5205 5630 6285
rect 5290 5175 5630 5205
rect 80 3320 145 5175
rect 1030 5135 1070 5175
rect 355 5125 1070 5135
rect 355 5105 1040 5125
rect 1060 5105 1070 5125
rect 355 5095 1070 5105
rect 355 4850 395 5095
rect 2615 5065 2655 5175
rect 1955 5025 2655 5065
rect 1955 4960 1995 5025
rect 3045 5005 3085 5175
rect 1955 4940 1965 4960
rect 1985 4940 1995 4960
rect 210 4820 550 4850
rect 1955 4845 1995 4940
rect 2390 4965 3085 5005
rect 2390 4845 2430 4965
rect 210 3740 240 4820
rect 520 3740 550 4820
rect 210 3710 550 3740
rect 1010 4820 1380 4845
rect 1010 3740 1040 4820
rect 1320 3740 1380 4820
rect 1010 3710 1380 3740
rect 1810 4820 2150 4845
rect 1810 3740 1840 4820
rect 2120 3740 2150 4820
rect 1810 3710 2150 3740
rect 2240 4820 2580 4845
rect 2240 3740 2270 4820
rect 2550 3740 2580 4820
rect 2240 3710 2580 3740
rect 3040 4820 3410 4845
rect 3040 3740 3070 4820
rect 3355 3740 3410 4820
rect 3040 3710 3410 3740
rect 1045 3520 1320 3710
rect 2385 3580 2425 3710
rect 2385 3560 2395 3580
rect 2415 3560 2425 3580
rect 2385 3550 2425 3560
rect 3045 3520 3410 3710
rect 3700 3610 3760 5175
rect 5440 5140 5480 5175
rect 3980 5125 5480 5140
rect 3980 5105 5450 5125
rect 5470 5105 5480 5125
rect 3980 5095 5480 5105
rect 3980 4850 4035 5095
rect 3835 4820 4175 4850
rect 3835 3740 3865 4820
rect 4145 3740 4175 4820
rect 3835 3710 4175 3740
rect 4245 4820 4615 4850
rect 4245 3740 4305 4820
rect 4585 3740 4615 4820
rect 4245 3710 4615 3740
rect 5075 4820 5705 4850
rect 5075 3740 5105 4820
rect 5385 4770 5705 4820
rect 5385 3740 5415 4770
rect 5075 3715 5415 3740
rect 5075 3710 5205 3715
rect 5275 3710 5415 3715
rect 3700 3555 3875 3610
rect 25 3250 145 3320
rect 80 1555 145 3250
rect 745 3465 1885 3520
rect 745 3185 770 3465
rect 1855 3185 1885 3465
rect 745 3130 1885 3185
rect 2580 3465 3720 3520
rect 2580 3185 2610 3465
rect 3690 3185 3720 3465
rect 2580 3135 3720 3185
rect 1045 2940 1320 3130
rect 2385 3090 2425 3100
rect 2385 3070 2395 3090
rect 2415 3070 2425 3090
rect 2385 2940 2425 3070
rect 3045 2940 3410 3135
rect 3815 3095 3875 3555
rect 4250 3520 4620 3710
rect 4080 3465 5220 3520
rect 4080 3185 4110 3465
rect 5190 3185 5220 3465
rect 4080 3135 5220 3185
rect 210 2910 550 2940
rect 210 1830 240 2910
rect 520 1830 550 2910
rect 210 1800 550 1830
rect 1010 2910 1380 2940
rect 1010 1830 1040 2910
rect 1325 1830 1380 2910
rect 1010 1805 1380 1830
rect 1810 2910 2150 2940
rect 1810 1830 1840 2910
rect 2120 1830 2150 2910
rect 1810 1800 2150 1830
rect 2240 2910 2580 2940
rect 2240 1830 2270 2910
rect 2550 1830 2580 2910
rect 2240 1800 2580 1830
rect 3040 2910 3410 2940
rect 3040 1830 3070 2910
rect 3350 1830 3410 2910
rect 3040 1800 3410 1830
rect 3700 3040 3875 3095
rect 350 1640 395 1800
rect 1955 1710 1995 1800
rect 1955 1690 1965 1710
rect 1985 1690 1995 1710
rect 1955 1640 1995 1690
rect 2390 1695 2430 1800
rect 2390 1660 3085 1695
rect 350 1625 1070 1640
rect 350 1605 1040 1625
rect 1060 1605 1070 1625
rect 350 1595 1070 1605
rect 1955 1600 2655 1640
rect 1030 1555 1070 1595
rect 2615 1555 2655 1600
rect 3045 1555 3085 1660
rect 3700 1555 3760 3040
rect 4250 2940 4620 3135
rect 5285 2940 5410 3710
rect 5665 3087 5705 3097
rect 5665 3027 5675 3087
rect 5695 3027 5705 3087
rect 5665 3017 5705 3027
rect 3835 2910 4175 2940
rect 3835 1830 3865 2910
rect 4145 1830 4175 2910
rect 3835 1800 4175 1830
rect 4245 2910 4620 2940
rect 4245 1830 4305 2910
rect 4585 2885 4620 2910
rect 5075 2910 5415 2940
rect 4585 1830 4615 2885
rect 4245 1800 4615 1830
rect 5075 1830 5105 2910
rect 5385 1830 5415 2910
rect 5075 1800 5415 1830
rect 3980 1640 4035 1800
rect 3980 1625 5480 1640
rect 3980 1605 5450 1625
rect 5470 1605 5480 1625
rect 3980 1595 5480 1605
rect 5440 1555 5480 1595
rect 80 1525 420 1555
rect 80 445 110 1525
rect 390 445 420 1525
rect 80 410 420 445
rect 880 1525 1220 1555
rect 880 445 910 1525
rect 1190 445 1220 1525
rect 880 415 1220 445
rect 1275 1525 2010 1555
rect 1275 445 1305 1525
rect 1590 445 1700 1525
rect 1985 445 2010 1525
rect 1275 415 2010 445
rect 2470 1525 2810 1555
rect 2470 445 2500 1525
rect 2780 445 2810 1525
rect 2470 415 2810 445
rect 2900 1525 3240 1555
rect 2900 445 2930 1525
rect 3210 445 3240 1525
rect 2900 415 3240 445
rect 3700 1525 4830 1555
rect 3700 445 3730 1525
rect 4015 445 4125 1525
rect 4410 445 4520 1525
rect 4805 445 4830 1525
rect 3700 415 4830 445
rect 5290 1525 5630 1555
rect 5290 445 5320 1525
rect 5600 445 5630 1525
rect 5290 415 5630 445
<< viali >>
rect 1300 5205 1305 6285
rect 1305 5205 1585 6285
rect 1695 5205 1700 6285
rect 1700 5205 1980 6285
rect 3730 5205 4010 6285
rect 4010 5205 4015 6285
rect 4120 5205 4125 6285
rect 4125 5205 4405 6285
rect 4520 5205 4800 6285
rect 4800 5205 4805 6285
rect 1040 3740 1320 4820
rect 3075 3740 3350 4820
rect 3350 3740 3355 4820
rect 4305 3740 4585 4820
rect 770 3185 775 3465
rect 775 3185 1850 3465
rect 2615 3185 3690 3465
rect 4110 3185 5185 3465
rect 1045 1830 1320 2910
rect 1320 1830 1325 2910
rect 3070 1830 3350 2910
rect 4305 1830 4585 2910
rect 1305 445 1585 1525
rect 1585 445 1590 1525
rect 1700 445 1980 1525
rect 1980 445 1985 1525
rect 3730 445 4010 1525
rect 4010 445 4015 1525
rect 4125 445 4405 1525
rect 4405 445 4410 1525
rect 4520 445 4800 1525
rect 4800 445 4805 1525
<< metal1 >>
rect 25 6285 5705 6350
rect 25 5205 1300 6285
rect 1585 5205 1695 6285
rect 1980 5205 3730 6285
rect 4015 5205 4120 6285
rect 4405 5205 4520 6285
rect 4805 5205 5705 6285
rect 25 5140 5705 5205
rect 25 4820 5705 4880
rect 25 3740 1040 4820
rect 1320 3740 3075 4820
rect 3355 3740 4305 4820
rect 4585 3740 5705 4820
rect 25 3465 5705 3740
rect 25 3185 770 3465
rect 1850 3185 2615 3465
rect 3690 3185 4110 3465
rect 5185 3185 5705 3465
rect 25 2910 5705 3185
rect 25 1830 1045 2910
rect 1325 1830 3070 2910
rect 3350 1830 4305 2910
rect 4585 1830 5705 2910
rect 25 1770 5705 1830
rect 25 1585 75 1590
rect 25 1525 5705 1585
rect 25 445 1305 1525
rect 1590 445 1700 1525
rect 1985 445 3730 1525
rect 4015 445 4125 1525
rect 4410 445 4520 1525
rect 4805 445 5705 1525
rect 25 385 5705 445
<< metal2 >>
rect 1969 6323 2160 6325
rect 1274 5176 2160 6323
rect 1969 1559 2160 5176
rect 1273 412 2160 1559
<< labels >>
flabel pmos 605 1795 900 2175 0 FreeSans 800 0 0 0 VG
flabel pmos 605 4475 900 4855 0 FreeSans 800 0 0 0 VG
rlabel locali 25 3285 25 3285 7 R
port 1 w
rlabel metal1 25 3365 25 3365 7 VP
port 2 w
rlabel locali 5705 4810 5705 4810 3 Ib
port 4 e
rlabel metal1 25 979 25 979 7 VN
port 3 w
rlabel locali 5705 3057 5705 3057 3 Vbn
port 5 e
<< end >>
