magic
tech sky130A
magscale 1 2
timestamp 1701147612
<< error_p >>
rect 39314 -9645 39315 -8348
rect 39314 -9646 39434 -9645
rect 39314 -11970 39315 -10106
<< nwell >>
rect -3820 -9470 2610 -6920
rect -3820 -9476 -3552 -9470
<< nmos >>
rect -3550 -11970 -3450 -9570
rect -3400 -11970 -3300 -9570
rect -3250 -11970 -3150 -9570
rect -3100 -11970 -3000 -9570
rect -2950 -11970 -2850 -9570
rect -2570 -11970 -2470 -9570
rect -2130 -11970 -2030 -9570
rect -1930 -11970 -1830 -9570
rect -1730 -11970 -1630 -9570
rect -1530 -11970 -1430 -9570
rect -1330 -11970 -1230 -9570
rect -1130 -11970 -1030 -9570
rect -770 -11970 -670 -9570
rect -400 -11970 -300 -9570
rect -40 -11970 60 -9570
rect 160 -11970 260 -9570
rect 360 -11970 460 -9570
rect 560 -11970 660 -9570
rect 760 -11970 860 -9570
rect 960 -11970 1060 -9570
rect 1400 -11970 1500 -9570
rect 1780 -11970 1880 -9570
rect 1930 -11970 2030 -9570
rect 2080 -11970 2180 -9570
rect 2230 -11970 2330 -9570
rect 2380 -11970 2480 -9570
<< pmos >>
rect -3460 -9370 -3360 -6970
rect -3260 -9370 -3160 -6970
rect -3060 -9370 -2960 -6970
rect -2860 -9370 -2760 -6970
rect -2660 -9370 -2560 -6970
rect -2460 -9370 -2360 -6970
rect -2100 -9370 -2000 -6970
rect -1950 -9370 -1850 -6970
rect -1800 -9370 -1700 -6970
rect -1650 -9370 -1550 -6970
rect -1500 -9370 -1400 -6970
rect -1130 -9370 -1030 -6970
rect -770 -9370 -670 -6970
rect -400 -9370 -300 -6970
rect -40 -9370 60 -6970
rect 330 -9370 430 -6970
rect 480 -9370 580 -6970
rect 630 -9370 730 -6970
rect 780 -9370 880 -6970
rect 930 -9370 1030 -6970
rect 1290 -9370 1390 -6970
rect 1490 -9370 1590 -6970
rect 1690 -9370 1790 -6970
rect 1890 -9370 1990 -6970
rect 2090 -9370 2190 -6970
rect 2290 -9370 2390 -6970
<< ndiff >>
rect -3650 -9600 -3550 -9570
rect -3650 -11940 -3620 -9600
rect -3580 -11940 -3550 -9600
rect -3650 -11970 -3550 -11940
rect -3450 -11970 -3400 -9570
rect -3300 -11970 -3250 -9570
rect -3150 -11970 -3100 -9570
rect -3000 -11970 -2950 -9570
rect -2850 -9600 -2750 -9570
rect -2670 -9600 -2570 -9570
rect -2850 -11940 -2820 -9600
rect -2780 -11940 -2750 -9600
rect -2670 -11940 -2640 -9600
rect -2600 -11940 -2570 -9600
rect -2850 -11970 -2750 -11940
rect -2670 -11970 -2570 -11940
rect -2470 -9600 -2370 -9570
rect -2470 -11940 -2440 -9600
rect -2400 -11940 -2370 -9600
rect -2470 -11970 -2370 -11940
rect -2220 -9600 -2130 -9570
rect -2220 -11940 -2200 -9600
rect -2160 -11940 -2130 -9600
rect -2220 -11970 -2130 -11940
rect -2030 -9600 -1930 -9570
rect -2030 -11940 -2000 -9600
rect -1960 -11940 -1930 -9600
rect -2030 -11970 -1930 -11940
rect -1830 -9600 -1730 -9570
rect -1830 -11940 -1800 -9600
rect -1760 -11940 -1730 -9600
rect -1830 -11970 -1730 -11940
rect -1630 -9600 -1530 -9570
rect -1630 -11940 -1600 -9600
rect -1560 -11940 -1530 -9600
rect -1630 -11970 -1530 -11940
rect -1430 -9600 -1330 -9570
rect -1430 -11940 -1400 -9600
rect -1360 -11940 -1330 -9600
rect -1430 -11970 -1330 -11940
rect -1230 -9600 -1130 -9570
rect -1230 -11940 -1200 -9600
rect -1160 -11940 -1130 -9600
rect -1230 -11970 -1130 -11940
rect -1030 -9600 -930 -9570
rect -1030 -11940 -1000 -9600
rect -960 -11940 -930 -9600
rect -1030 -11970 -930 -11940
rect -870 -9600 -770 -9570
rect -870 -11940 -840 -9600
rect -800 -11940 -770 -9600
rect -870 -11970 -770 -11940
rect -670 -9600 -580 -9570
rect -500 -9600 -400 -9570
rect -670 -11940 -650 -9600
rect -610 -11940 -580 -9600
rect -500 -11940 -470 -9600
rect -430 -11940 -400 -9600
rect -670 -11970 -580 -11940
rect -500 -11970 -400 -11940
rect -300 -9600 -200 -9570
rect -300 -11940 -270 -9600
rect -230 -11940 -200 -9600
rect -300 -11970 -200 -11940
rect -140 -9600 -40 -9570
rect -140 -11940 -110 -9600
rect -70 -11940 -40 -9600
rect -140 -11970 -40 -11940
rect 60 -9600 160 -9570
rect 60 -11940 90 -9600
rect 130 -11940 160 -9600
rect 60 -11970 160 -11940
rect 260 -9600 360 -9570
rect 260 -11940 290 -9600
rect 330 -11940 360 -9600
rect 260 -11970 360 -11940
rect 460 -9600 560 -9570
rect 460 -11940 490 -9600
rect 530 -11940 560 -9600
rect 460 -11970 560 -11940
rect 660 -9600 760 -9570
rect 660 -11940 690 -9600
rect 730 -11940 760 -9600
rect 660 -11970 760 -11940
rect 860 -9600 960 -9570
rect 860 -11940 890 -9600
rect 930 -11940 960 -9600
rect 860 -11970 960 -11940
rect 1060 -9600 1150 -9570
rect 1060 -11940 1090 -9600
rect 1130 -11940 1150 -9600
rect 1060 -11970 1150 -11940
rect 1300 -9600 1400 -9570
rect 1300 -11940 1330 -9600
rect 1370 -11940 1400 -9600
rect 1300 -11970 1400 -11940
rect 1500 -9600 1600 -9570
rect 1680 -9600 1780 -9570
rect 1500 -11940 1530 -9600
rect 1570 -11940 1600 -9600
rect 1680 -11940 1710 -9600
rect 1750 -11940 1780 -9600
rect 1500 -11970 1600 -11940
rect 1680 -11970 1780 -11940
rect 1880 -11970 1930 -9570
rect 2030 -11970 2080 -9570
rect 2180 -11970 2230 -9570
rect 2330 -11970 2380 -9570
rect 2480 -9600 2580 -9570
rect 2480 -11940 2510 -9600
rect 2550 -11940 2580 -9600
rect 2480 -11970 2580 -11940
<< pdiff >>
rect -3550 -7000 -3460 -6970
rect -3550 -9340 -3530 -7000
rect -3490 -9340 -3460 -7000
rect -3550 -9370 -3460 -9340
rect -3360 -7000 -3260 -6970
rect -3360 -9340 -3330 -7000
rect -3290 -9340 -3260 -7000
rect -3360 -9370 -3260 -9340
rect -3160 -7000 -3060 -6970
rect -3160 -9340 -3130 -7000
rect -3090 -9340 -3060 -7000
rect -3160 -9370 -3060 -9340
rect -2960 -7000 -2860 -6970
rect -2960 -9340 -2930 -7000
rect -2890 -9340 -2860 -7000
rect -2960 -9370 -2860 -9340
rect -2760 -7000 -2660 -6970
rect -2760 -9340 -2730 -7000
rect -2690 -9340 -2660 -7000
rect -2760 -9370 -2660 -9340
rect -2560 -7000 -2460 -6970
rect -2560 -9340 -2530 -7000
rect -2490 -9340 -2460 -7000
rect -2560 -9370 -2460 -9340
rect -2360 -7000 -2260 -6970
rect -2360 -9340 -2330 -7000
rect -2290 -9340 -2260 -7000
rect -2360 -9370 -2260 -9340
rect -2200 -7000 -2100 -6970
rect -2200 -9340 -2170 -7000
rect -2130 -9340 -2100 -7000
rect -2200 -9370 -2100 -9340
rect -2000 -9370 -1950 -6970
rect -1850 -9370 -1800 -6970
rect -1700 -9370 -1650 -6970
rect -1550 -9370 -1500 -6970
rect -1400 -7000 -1300 -6970
rect -1220 -7000 -1130 -6970
rect -1400 -9340 -1370 -7000
rect -1330 -9340 -1300 -7000
rect -1220 -9340 -1200 -7000
rect -1160 -9340 -1130 -7000
rect -1400 -9370 -1300 -9340
rect -1220 -9370 -1130 -9340
rect -1030 -7000 -930 -6970
rect -1030 -9340 -1000 -7000
rect -960 -9340 -930 -7000
rect -1030 -9370 -930 -9340
rect -870 -7000 -770 -6970
rect -870 -9340 -840 -7000
rect -800 -9340 -770 -7000
rect -870 -9370 -770 -9340
rect -670 -7000 -580 -6970
rect -500 -7000 -400 -6970
rect -670 -9340 -640 -7000
rect -600 -9340 -580 -7000
rect -500 -9340 -470 -7000
rect -430 -9340 -400 -7000
rect -670 -9370 -580 -9340
rect -500 -9370 -400 -9340
rect -300 -7000 -200 -6970
rect -300 -9340 -270 -7000
rect -230 -9340 -200 -7000
rect -300 -9370 -200 -9340
rect -140 -7000 -40 -6970
rect -140 -9340 -110 -7000
rect -70 -9340 -40 -7000
rect -140 -9370 -40 -9340
rect 60 -7000 150 -6970
rect 230 -7000 330 -6970
rect 60 -9340 90 -7000
rect 130 -9340 150 -7000
rect 230 -9340 260 -7000
rect 300 -9340 330 -7000
rect 60 -9370 150 -9340
rect 230 -9370 330 -9340
rect 430 -9370 480 -6970
rect 580 -9370 630 -6970
rect 730 -9370 780 -6970
rect 880 -9370 930 -6970
rect 1030 -7000 1130 -6970
rect 1030 -9340 1060 -7000
rect 1100 -9340 1130 -7000
rect 1030 -9370 1130 -9340
rect 1190 -7000 1290 -6970
rect 1190 -9340 1220 -7000
rect 1260 -9340 1290 -7000
rect 1190 -9370 1290 -9340
rect 1390 -7000 1490 -6970
rect 1390 -9340 1420 -7000
rect 1460 -9340 1490 -7000
rect 1390 -9370 1490 -9340
rect 1590 -7000 1690 -6970
rect 1590 -9340 1620 -7000
rect 1660 -9340 1690 -7000
rect 1590 -9370 1690 -9340
rect 1790 -7000 1890 -6970
rect 1790 -9340 1820 -7000
rect 1860 -9340 1890 -7000
rect 1790 -9370 1890 -9340
rect 1990 -7000 2090 -6970
rect 1990 -9340 2020 -7000
rect 2060 -9340 2090 -7000
rect 1990 -9370 2090 -9340
rect 2190 -7000 2290 -6970
rect 2190 -9340 2220 -7000
rect 2260 -9340 2290 -7000
rect 2190 -9370 2290 -9340
rect 2390 -7000 2480 -6970
rect 2390 -9340 2420 -7000
rect 2460 -9340 2480 -7000
rect 2390 -9370 2480 -9340
<< ndiffc >>
rect -3620 -11940 -3580 -9600
rect -2820 -11940 -2780 -9600
rect -2640 -11940 -2600 -9600
rect -2440 -11940 -2400 -9600
rect -2200 -11940 -2160 -9600
rect -2000 -11940 -1960 -9600
rect -1800 -11940 -1760 -9600
rect -1600 -11940 -1560 -9600
rect -1400 -11940 -1360 -9600
rect -1200 -11940 -1160 -9600
rect -1000 -11940 -960 -9600
rect -840 -11940 -800 -9600
rect -650 -11940 -610 -9600
rect -470 -11940 -430 -9600
rect -270 -11940 -230 -9600
rect -110 -11940 -70 -9600
rect 90 -11940 130 -9600
rect 290 -11940 330 -9600
rect 490 -11940 530 -9600
rect 690 -11940 730 -9600
rect 890 -11940 930 -9600
rect 1090 -11940 1130 -9600
rect 1330 -11940 1370 -9600
rect 1530 -11940 1570 -9600
rect 1710 -11940 1750 -9600
rect 2510 -11940 2550 -9600
<< pdiffc >>
rect -3530 -9340 -3490 -7000
rect -3330 -9340 -3290 -7000
rect -3130 -9340 -3090 -7000
rect -2930 -9340 -2890 -7000
rect -2730 -9340 -2690 -7000
rect -2530 -9340 -2490 -7000
rect -2330 -9340 -2290 -7000
rect -2170 -9340 -2130 -7000
rect -1370 -9340 -1330 -7000
rect -1200 -9340 -1160 -7000
rect -1000 -9340 -960 -7000
rect -840 -9340 -800 -7000
rect -640 -9340 -600 -7000
rect -470 -9340 -430 -7000
rect -270 -9340 -230 -7000
rect -110 -9340 -70 -7000
rect 90 -9340 130 -7000
rect 260 -9340 300 -7000
rect 1060 -9340 1100 -7000
rect 1220 -9340 1260 -7000
rect 1420 -9340 1460 -7000
rect 1620 -9340 1660 -7000
rect 1820 -9340 1860 -7000
rect 2020 -9340 2060 -7000
rect 2220 -9340 2260 -7000
rect 2420 -9340 2460 -7000
<< psubdiff >>
rect -2750 -9600 -2670 -9570
rect -2750 -11940 -2730 -9600
rect -2690 -11940 -2670 -9600
rect -2750 -11970 -2670 -11940
rect -2310 -9600 -2220 -9570
rect -2310 -11940 -2280 -9600
rect -2240 -11940 -2220 -9600
rect -2310 -11970 -2220 -11940
rect -580 -9600 -500 -9570
rect -580 -11940 -560 -9600
rect -520 -11940 -500 -9600
rect -580 -11970 -500 -11940
rect 1150 -9600 1240 -9570
rect 1150 -11940 1170 -9600
rect 1210 -11940 1240 -9600
rect 1150 -11970 1240 -11940
rect 1600 -9600 1680 -9570
rect 1600 -11940 1620 -9600
rect 1660 -11940 1680 -9600
rect 1600 -11970 1680 -11940
<< nsubdiff >>
rect -3640 -7000 -3550 -6970
rect -3640 -9340 -3610 -7000
rect -3570 -9340 -3550 -7000
rect -3640 -9370 -3550 -9340
rect -1300 -7000 -1220 -6970
rect -1300 -9340 -1280 -7000
rect -1240 -9340 -1220 -7000
rect -1300 -9370 -1220 -9340
rect -580 -7000 -500 -6970
rect -580 -9340 -560 -7000
rect -520 -9340 -500 -7000
rect -580 -9370 -500 -9340
rect 150 -7000 230 -6970
rect 150 -9340 170 -7000
rect 210 -9340 230 -7000
rect 150 -9370 230 -9340
rect 2480 -7000 2570 -6970
rect 2480 -9340 2500 -7000
rect 2540 -9340 2570 -7000
rect 2480 -9370 2570 -9340
<< psubdiffcont >>
rect -2730 -11940 -2690 -9600
rect -2280 -11940 -2240 -9600
rect -560 -11940 -520 -9600
rect 1170 -11940 1210 -9600
rect 1620 -11940 1660 -9600
<< nsubdiffcont >>
rect -3610 -9340 -3570 -7000
rect -1280 -9340 -1240 -7000
rect -560 -9340 -520 -7000
rect 170 -9340 210 -7000
rect 2500 -9340 2540 -7000
<< poly >>
rect 35896 -3938 36702 -3936
rect 35232 -3970 36702 -3938
rect 35232 -4168 36326 -3970
rect 36668 -4168 36702 -3970
rect 35232 -4204 36702 -4168
rect -1130 -6650 -1030 -6640
rect -1130 -6690 -1100 -6650
rect -1060 -6690 -1030 -6650
rect -1130 -6860 -1030 -6690
rect -2100 -6890 -1030 -6860
rect -3460 -6970 -3360 -6940
rect -3260 -6970 -3160 -6940
rect -3060 -6970 -2960 -6940
rect -2860 -6970 -2760 -6940
rect -2660 -6970 -2560 -6940
rect -2460 -6970 -2360 -6940
rect -2100 -6970 -2000 -6890
rect -1950 -6970 -1850 -6890
rect -1800 -6970 -1700 -6890
rect -1650 -6970 -1550 -6890
rect -1500 -6970 -1400 -6890
rect -1130 -6970 -1030 -6890
rect -770 -6650 -670 -6640
rect -770 -6690 -740 -6650
rect -700 -6690 -670 -6650
rect -770 -6970 -670 -6690
rect -400 -6650 -300 -6640
rect -400 -6690 -370 -6650
rect -330 -6690 -300 -6650
rect -400 -6970 -300 -6690
rect -40 -6650 60 -6640
rect -40 -6690 -10 -6650
rect 30 -6690 60 -6650
rect -40 -6860 60 -6690
rect -40 -6890 1030 -6860
rect -40 -6970 60 -6890
rect 330 -6970 430 -6890
rect 480 -6970 580 -6890
rect 630 -6970 730 -6890
rect 780 -6970 880 -6890
rect 930 -6970 1030 -6890
rect 1290 -6970 1390 -6940
rect 1490 -6970 1590 -6940
rect 1690 -6970 1790 -6940
rect 1890 -6970 1990 -6940
rect 2090 -6970 2190 -6940
rect 2290 -6970 2390 -6940
rect -3650 -9420 -3550 -9410
rect -3650 -9460 -3620 -9420
rect -3580 -9440 -3550 -9420
rect -3460 -9440 -3360 -9370
rect -3260 -9410 -3160 -9370
rect -3060 -9410 -2960 -9370
rect -3260 -9420 -2960 -9410
rect -3260 -9440 -3130 -9420
rect -3580 -9460 -3130 -9440
rect -3090 -9440 -2960 -9420
rect -2860 -9410 -2760 -9370
rect -2660 -9410 -2560 -9370
rect -2860 -9420 -2560 -9410
rect -2860 -9440 -2730 -9420
rect -3090 -9460 -2730 -9440
rect -2690 -9460 -2560 -9420
rect -3650 -9470 -2560 -9460
rect -2460 -9410 -2360 -9370
rect -2100 -9400 -2000 -9370
rect -1950 -9400 -1850 -9370
rect -1800 -9400 -1700 -9370
rect -1650 -9400 -1550 -9370
rect -1500 -9400 -1400 -9370
rect -1130 -9400 -1030 -9370
rect -770 -9400 -670 -9370
rect -400 -9400 -300 -9370
rect -40 -9400 60 -9370
rect 330 -9400 430 -9370
rect 480 -9400 580 -9370
rect 630 -9400 730 -9370
rect 780 -9400 880 -9370
rect 930 -9400 1030 -9370
rect 1290 -9410 1390 -9370
rect -2460 -9420 -2260 -9410
rect -2460 -9460 -2330 -9420
rect -2290 -9460 -2260 -9420
rect 1190 -9420 1390 -9410
rect -2460 -9470 -2260 -9460
rect -2200 -9460 -2030 -9450
rect -2200 -9500 -2170 -9460
rect -2130 -9500 -2030 -9460
rect -2200 -9510 -2030 -9500
rect -3550 -9570 -3450 -9540
rect -3400 -9570 -3300 -9540
rect -3250 -9570 -3150 -9540
rect -3100 -9570 -3000 -9540
rect -2950 -9570 -2850 -9540
rect -2570 -9570 -2470 -9540
rect -2130 -9570 -2030 -9510
rect 960 -9460 1130 -9450
rect 960 -9500 1060 -9460
rect 1100 -9500 1130 -9460
rect 1190 -9460 1220 -9420
rect 1260 -9460 1390 -9420
rect 1190 -9470 1390 -9460
rect 1490 -9410 1590 -9370
rect 1690 -9410 1790 -9370
rect 1490 -9420 1790 -9410
rect 1490 -9460 1620 -9420
rect 1660 -9440 1790 -9420
rect 1890 -9410 1990 -9370
rect 2090 -9410 2190 -9370
rect 1890 -9420 2190 -9410
rect 1890 -9440 2020 -9420
rect 1660 -9460 2020 -9440
rect 2060 -9440 2190 -9420
rect 2290 -9440 2390 -9370
rect 2480 -9420 2580 -9410
rect 2480 -9440 2510 -9420
rect 2060 -9460 2510 -9440
rect 2550 -9460 2580 -9420
rect 1490 -9470 2580 -9460
rect 960 -9510 1130 -9500
rect -1930 -9570 -1830 -9540
rect -1730 -9570 -1630 -9540
rect -1530 -9570 -1430 -9540
rect -1330 -9570 -1230 -9540
rect -1130 -9570 -1030 -9540
rect -770 -9570 -670 -9540
rect -400 -9570 -300 -9540
rect -40 -9570 60 -9540
rect 160 -9570 260 -9540
rect 360 -9570 460 -9540
rect 560 -9570 660 -9540
rect 760 -9570 860 -9540
rect 960 -9570 1060 -9510
rect 1400 -9570 1500 -9540
rect 1780 -9570 1880 -9540
rect 1930 -9570 2030 -9540
rect 2080 -9570 2180 -9540
rect 2230 -9570 2330 -9540
rect 2380 -9570 2480 -9540
rect -3550 -12030 -3450 -11970
rect -3400 -12030 -3300 -11970
rect -3250 -12030 -3150 -11970
rect -3100 -12030 -3000 -11970
rect -2950 -12030 -2850 -11970
rect -2570 -12030 -2470 -11970
rect -3550 -12060 -2470 -12030
rect -2570 -12220 -2470 -12060
rect -2130 -12040 -2030 -11970
rect -1930 -12010 -1830 -11970
rect -1730 -12010 -1630 -11970
rect -1930 -12020 -1630 -12010
rect -1930 -12040 -1800 -12020
rect -2130 -12060 -1800 -12040
rect -1760 -12040 -1630 -12020
rect -1530 -12010 -1430 -11970
rect -1330 -12010 -1230 -11970
rect -1530 -12020 -1230 -12010
rect -1530 -12040 -1400 -12020
rect -1760 -12060 -1400 -12040
rect -1360 -12060 -1230 -12020
rect -2130 -12070 -1230 -12060
rect -1130 -12000 -1030 -11970
rect -1130 -12010 -930 -12000
rect -1130 -12050 -1000 -12010
rect -960 -12050 -930 -12010
rect -1130 -12060 -930 -12050
rect -770 -12010 -670 -11970
rect -770 -12050 -740 -12010
rect -700 -12050 -670 -12010
rect -770 -12060 -670 -12050
rect -400 -12010 -300 -11970
rect -40 -12000 60 -11970
rect -400 -12050 -370 -12010
rect -330 -12050 -300 -12010
rect -400 -12060 -300 -12050
rect -140 -12010 60 -12000
rect -140 -12050 -110 -12010
rect -70 -12050 60 -12010
rect -140 -12060 60 -12050
rect -1130 -12110 -1030 -12060
rect -40 -12110 60 -12060
rect 160 -12010 260 -11970
rect 360 -12010 460 -11970
rect 160 -12020 460 -12010
rect 160 -12060 290 -12020
rect 330 -12040 460 -12020
rect 560 -12010 660 -11970
rect 760 -12010 860 -11970
rect 560 -12020 860 -12010
rect 560 -12040 690 -12020
rect 330 -12060 690 -12040
rect 730 -12040 860 -12020
rect 960 -12040 1060 -11970
rect 730 -12060 1060 -12040
rect 160 -12070 1060 -12060
rect 1400 -12030 1500 -11970
rect 1780 -12030 1880 -11970
rect 1930 -12030 2030 -11970
rect 2080 -12030 2180 -11970
rect 2230 -12030 2330 -11970
rect 2380 -12030 2480 -11970
rect 1400 -12060 2480 -12030
rect -1130 -12160 60 -12110
rect -2570 -12260 -2540 -12220
rect -2500 -12260 -2470 -12220
rect -2570 -12270 -2470 -12260
rect 1400 -12220 1500 -12060
rect 1400 -12260 1430 -12220
rect 1470 -12260 1500 -12220
rect 1400 -12270 1500 -12260
<< polycont >>
rect 36326 -4168 36668 -3970
rect -1100 -6690 -1060 -6650
rect -740 -6690 -700 -6650
rect -370 -6690 -330 -6650
rect -10 -6690 30 -6650
rect -3620 -9460 -3580 -9420
rect -3130 -9460 -3090 -9420
rect -2730 -9460 -2690 -9420
rect -2330 -9460 -2290 -9420
rect -2170 -9500 -2130 -9460
rect 1060 -9500 1100 -9460
rect 1220 -9460 1260 -9420
rect 1620 -9460 1660 -9420
rect 2020 -9460 2060 -9420
rect 2510 -9460 2550 -9420
rect -1800 -12060 -1760 -12020
rect -1400 -12060 -1360 -12020
rect -1000 -12050 -960 -12010
rect -740 -12050 -700 -12010
rect -370 -12050 -330 -12010
rect -110 -12050 -70 -12010
rect 290 -12060 330 -12020
rect 690 -12060 730 -12020
rect -2540 -12260 -2500 -12220
rect 1430 -12260 1470 -12220
rect 4100 -15410 4240 -15250
rect 4100 -20770 4340 -20630
<< locali >>
rect 30610 -1166 31032 -1152
rect 30610 -1356 30626 -1166
rect 31016 -1356 31032 -1166
rect 30610 -1370 31032 -1356
rect 30682 -1432 31032 -1416
rect 30682 -1468 30692 -1432
rect 30958 -1468 31032 -1432
rect 30682 -1472 31032 -1468
rect 30682 -1476 30968 -1472
rect -3820 -2930 -2900 -2830
rect -3820 -3110 -3640 -2930
rect -3080 -3110 -2900 -2930
rect -3820 -3210 -2900 -3110
rect 36288 -3970 36702 -3936
rect 36288 -4168 36326 -3970
rect 36668 -4168 36702 -3970
rect 36288 -4204 36702 -4168
rect -3820 -6650 2750 -6640
rect -3820 -6690 -1100 -6650
rect -1060 -6690 -740 -6650
rect -700 -6690 -370 -6650
rect -330 -6690 -10 -6650
rect 30 -6690 2660 -6650
rect 2740 -6690 2750 -6650
rect -3820 -6700 2750 -6690
rect 30882 -6732 31032 -6718
rect -2350 -6768 4722 -6760
rect -2350 -6812 3974 -6768
rect 4710 -6812 4722 -6768
rect -2350 -6820 4722 -6812
rect -3350 -6940 -2460 -6870
rect -3630 -6980 -3550 -6960
rect -3630 -7000 -3470 -6980
rect -3630 -9340 -3610 -7000
rect -3570 -9340 -3530 -7000
rect -3490 -9340 -3470 -7000
rect -3630 -9360 -3470 -9340
rect -3350 -7000 -3270 -6940
rect -3350 -9340 -3330 -7000
rect -3290 -9340 -3270 -7000
rect -3350 -9360 -3270 -9340
rect -3150 -7000 -3070 -6980
rect -3150 -9340 -3130 -7000
rect -3090 -9340 -3070 -7000
rect -3150 -9410 -3070 -9340
rect -2950 -7000 -2870 -6940
rect -2950 -9340 -2930 -7000
rect -2890 -9340 -2870 -7000
rect -2950 -9360 -2870 -9340
rect -2750 -7000 -2670 -6980
rect -2750 -9340 -2730 -7000
rect -2690 -9340 -2670 -7000
rect -2750 -9410 -2670 -9340
rect -2550 -7000 -2460 -6940
rect -2550 -9340 -2530 -7000
rect -2490 -9340 -2460 -7000
rect -2550 -9360 -2460 -9340
rect -2350 -7000 -2270 -6820
rect -2350 -9340 -2330 -7000
rect -2290 -9340 -2270 -7000
rect -2350 -9410 -2270 -9340
rect -2190 -7000 -2110 -6980
rect -2190 -9340 -2170 -7000
rect -2130 -9340 -2110 -7000
rect -3650 -9420 -3550 -9410
rect -3650 -9460 -3620 -9420
rect -3580 -9460 -3550 -9420
rect -3650 -9470 -3550 -9460
rect -3160 -9420 -3060 -9410
rect -3160 -9460 -3130 -9420
rect -3090 -9460 -3060 -9420
rect -3160 -9470 -3060 -9460
rect -2760 -9420 -2660 -9410
rect -2760 -9460 -2730 -9420
rect -2690 -9460 -2660 -9420
rect -2760 -9470 -2660 -9460
rect -2460 -9420 -2260 -9410
rect -2460 -9460 -2330 -9420
rect -2290 -9460 -2260 -9420
rect -2190 -9450 -2110 -9340
rect -1390 -7000 -1140 -6980
rect -1390 -9340 -1370 -7000
rect -1330 -9340 -1280 -7000
rect -1240 -9340 -1200 -7000
rect -1160 -9340 -1140 -7000
rect -1390 -9360 -1140 -9340
rect -1020 -7000 -940 -6980
rect -1020 -9340 -1000 -7000
rect -960 -9340 -940 -7000
rect -2460 -9470 -2260 -9460
rect -2200 -9460 -2100 -9450
rect -3640 -9600 -3560 -9470
rect -3640 -11940 -3620 -9600
rect -3580 -11940 -3560 -9600
rect -3640 -11960 -3560 -11940
rect -2840 -9600 -2580 -9580
rect -2840 -11940 -2820 -9600
rect -2770 -11940 -2730 -9600
rect -2690 -11940 -2650 -9600
rect -2600 -11940 -2580 -9600
rect -2840 -11960 -2580 -11940
rect -2460 -9600 -2380 -9470
rect -2200 -9500 -2170 -9460
rect -2130 -9500 -2100 -9460
rect -2200 -9510 -2100 -9500
rect -2020 -9540 -1130 -9470
rect -2460 -11940 -2440 -9600
rect -2400 -11940 -2380 -9600
rect -2460 -11960 -2380 -11940
rect -2300 -9600 -2140 -9580
rect -2300 -11940 -2280 -9600
rect -2240 -11940 -2200 -9600
rect -2160 -11940 -2140 -9600
rect -2300 -11960 -2140 -11940
rect -2020 -9600 -1940 -9540
rect -2020 -11940 -2000 -9600
rect -1960 -11940 -1940 -9600
rect -2020 -11960 -1940 -11940
rect -1820 -9600 -1740 -9580
rect -1820 -11940 -1800 -9600
rect -1760 -11940 -1740 -9600
rect -1820 -12010 -1740 -11940
rect -1620 -9600 -1540 -9540
rect -1620 -11940 -1600 -9600
rect -1560 -11940 -1540 -9600
rect -1620 -11960 -1540 -11940
rect -1420 -9600 -1340 -9580
rect -1420 -11940 -1400 -9600
rect -1360 -11940 -1340 -9600
rect -1420 -12010 -1340 -11940
rect -1220 -9600 -1130 -9540
rect -1220 -11940 -1200 -9600
rect -1160 -11940 -1130 -9600
rect -1220 -11960 -1130 -11940
rect -1020 -9600 -940 -9340
rect -1020 -11940 -1000 -9600
rect -960 -11940 -940 -9600
rect -1020 -12000 -940 -11940
rect -860 -7000 -780 -6980
rect -860 -9340 -840 -7000
rect -800 -9340 -780 -7000
rect -860 -9600 -780 -9340
rect -670 -7000 -410 -6980
rect -670 -9340 -640 -7000
rect -600 -9340 -560 -7000
rect -520 -9340 -470 -7000
rect -430 -9340 -410 -7000
rect -670 -9360 -410 -9340
rect -290 -7000 -210 -6980
rect -290 -9340 -270 -7000
rect -230 -9340 -210 -7000
rect -860 -11940 -840 -9600
rect -800 -11940 -780 -9600
rect -860 -12000 -780 -11940
rect -670 -9600 -410 -9580
rect -670 -11940 -650 -9600
rect -600 -11940 -560 -9600
rect -520 -11940 -480 -9600
rect -430 -11940 -410 -9600
rect -670 -11960 -410 -11940
rect -290 -9600 -210 -9340
rect -290 -11940 -270 -9600
rect -230 -11940 -210 -9600
rect -290 -12000 -210 -11940
rect -130 -7000 -50 -6980
rect -130 -9340 -110 -7000
rect -70 -9340 -50 -7000
rect -130 -9600 -50 -9340
rect 70 -7000 320 -6980
rect 70 -9340 90 -7000
rect 130 -9340 170 -7000
rect 210 -9340 260 -7000
rect 300 -9340 320 -7000
rect 70 -9360 320 -9340
rect 1040 -7000 1120 -6980
rect 1040 -9340 1060 -7000
rect 1100 -9340 1120 -7000
rect 1040 -9450 1120 -9340
rect 1200 -7000 1280 -6820
rect 30882 -6852 30896 -6732
rect 31016 -6852 31032 -6732
rect 30882 -6866 31032 -6852
rect 1200 -9340 1220 -7000
rect 1260 -9340 1280 -7000
rect 1200 -9410 1280 -9340
rect 1390 -6940 2280 -6870
rect 1390 -7000 1480 -6940
rect 1390 -9340 1420 -7000
rect 1460 -9340 1480 -7000
rect 1390 -9360 1480 -9340
rect 1600 -7000 1680 -6980
rect 1600 -9340 1620 -7000
rect 1660 -9340 1680 -7000
rect 1600 -9410 1680 -9340
rect 1800 -7000 1880 -6940
rect 1800 -9340 1820 -7000
rect 1860 -9340 1880 -7000
rect 1800 -9360 1880 -9340
rect 2000 -7000 2080 -6980
rect 2000 -9340 2020 -7000
rect 2060 -9340 2080 -7000
rect 2000 -9410 2080 -9340
rect 2200 -7000 2280 -6940
rect 2480 -6980 2560 -6960
rect 2200 -9340 2220 -7000
rect 2260 -9340 2280 -7000
rect 2200 -9360 2280 -9340
rect 2400 -7000 2560 -6980
rect 2400 -9340 2420 -7000
rect 2460 -9340 2500 -7000
rect 2540 -9340 2560 -7000
rect 2400 -9360 2560 -9340
rect 1190 -9420 1390 -9410
rect 1030 -9460 1130 -9450
rect -130 -11940 -110 -9600
rect -70 -11940 -50 -9600
rect -130 -12000 -50 -11940
rect 60 -9540 950 -9470
rect 1030 -9500 1060 -9460
rect 1100 -9500 1130 -9460
rect 1190 -9460 1220 -9420
rect 1260 -9460 1390 -9420
rect 1190 -9470 1390 -9460
rect 1590 -9420 1690 -9410
rect 1590 -9460 1620 -9420
rect 1660 -9460 1690 -9420
rect 1590 -9470 1690 -9460
rect 1990 -9420 2090 -9410
rect 1990 -9460 2020 -9420
rect 2060 -9460 2090 -9420
rect 1990 -9470 2090 -9460
rect 2480 -9420 2580 -9410
rect 2480 -9460 2510 -9420
rect 2550 -9460 2580 -9420
rect 2480 -9470 2580 -9460
rect 1030 -9510 1130 -9500
rect 60 -9600 150 -9540
rect 60 -11940 90 -9600
rect 130 -11940 150 -9600
rect 60 -11960 150 -11940
rect 270 -9600 350 -9580
rect 270 -11940 290 -9600
rect 330 -11940 350 -9600
rect -1030 -12010 -930 -12000
rect -1830 -12020 -1730 -12010
rect -1830 -12060 -1800 -12020
rect -1760 -12060 -1730 -12020
rect -1830 -12070 -1730 -12060
rect -1430 -12020 -1330 -12010
rect -1430 -12060 -1400 -12020
rect -1360 -12060 -1330 -12020
rect -1030 -12050 -1000 -12010
rect -960 -12050 -930 -12010
rect -1030 -12060 -930 -12050
rect -860 -12010 -670 -12000
rect -860 -12050 -740 -12010
rect -700 -12050 -670 -12010
rect -860 -12060 -670 -12050
rect -1430 -12070 -1330 -12060
rect -2570 -12220 -2470 -12210
rect -770 -12220 -670 -12060
rect -400 -12010 -210 -12000
rect -400 -12050 -370 -12010
rect -330 -12050 -210 -12010
rect -400 -12060 -210 -12050
rect -140 -12010 -40 -12000
rect 270 -12010 350 -11940
rect 470 -9600 550 -9540
rect 470 -11940 490 -9600
rect 530 -11940 550 -9600
rect 470 -11960 550 -11940
rect 670 -9600 750 -9580
rect 670 -11940 690 -9600
rect 730 -11940 750 -9600
rect 670 -12010 750 -11940
rect 870 -9600 950 -9540
rect 870 -11940 890 -9600
rect 930 -11940 950 -9600
rect 870 -11960 950 -11940
rect 1070 -9600 1230 -9580
rect 1070 -11940 1090 -9600
rect 1130 -11940 1170 -9600
rect 1210 -11940 1230 -9600
rect 1070 -11960 1230 -11940
rect 1310 -9600 1390 -9470
rect 1310 -11940 1330 -9600
rect 1370 -11940 1390 -9600
rect 1310 -11960 1390 -11940
rect 1510 -9600 1770 -9580
rect 1510 -11940 1530 -9600
rect 1580 -11940 1620 -9600
rect 1660 -11940 1700 -9600
rect 1750 -11940 1770 -9600
rect 1510 -11960 1770 -11940
rect 2490 -9600 2570 -9470
rect 2490 -11940 2510 -9600
rect 2550 -11940 2570 -9600
rect 35832 -9686 36794 -7366
rect 36288 -9812 36794 -9786
rect 36288 -9944 36318 -9812
rect 36662 -9944 36794 -9812
rect 36288 -9966 36794 -9944
rect 2490 -11960 2570 -11940
rect -140 -12050 -110 -12010
rect -70 -12050 -40 -12010
rect -400 -12220 -300 -12060
rect -140 -12120 -40 -12050
rect 260 -12020 360 -12010
rect 260 -12060 290 -12020
rect 330 -12060 360 -12020
rect 260 -12070 360 -12060
rect 660 -12020 760 -12010
rect 660 -12060 690 -12020
rect 730 -12060 760 -12020
rect 660 -12070 760 -12060
rect -140 -12170 2922 -12120
rect 1400 -12220 1500 -12210
rect -2570 -12260 -2540 -12220
rect -2500 -12260 1430 -12220
rect 1470 -12260 1500 -12220
rect -2570 -12270 1500 -12260
rect 2790 -12380 2922 -12170
rect 2790 -12458 2924 -12380
rect 2582 -12486 2924 -12458
rect 29864 -12468 31032 -12122
rect 35832 -12386 36794 -10066
rect 2582 -12816 2608 -12486
rect 2892 -12816 2924 -12486
rect 2582 -12844 2924 -12816
rect 2790 -12846 2924 -12844
rect 29866 -14764 30414 -12468
rect 29280 -14786 30414 -14764
rect 29280 -15148 29302 -14786
rect 29806 -15148 30414 -14786
rect 29280 -15172 30414 -15148
rect 30570 -15018 31032 -15000
rect 30570 -15158 30842 -15018
rect 31018 -15158 31032 -15018
rect 4060 -15250 4280 -15210
rect 4060 -15410 4100 -15250
rect 4240 -15410 4280 -15250
rect 4060 -15430 4280 -15410
rect 30570 -15482 31032 -15158
rect 2220 -15590 4580 -15530
rect 2220 -17790 2300 -15590
rect 2660 -17790 4140 -15590
rect 4500 -17790 4580 -15590
rect 30568 -15616 31032 -15482
rect 30568 -16066 31030 -15616
rect 30566 -16098 31030 -16066
rect 30566 -16530 31028 -16098
rect 30564 -16682 31028 -16530
rect 30564 -16950 31026 -16682
rect 2220 -18230 4580 -17790
rect 30562 -17146 31026 -16950
rect 30562 -18114 31024 -17146
rect 2220 -18250 4140 -18230
rect 2220 -20450 2300 -18250
rect 2660 -20430 4140 -18250
rect 4500 -20430 4580 -18230
rect 30560 -18180 31024 -18114
rect 30560 -18560 31022 -18180
rect 2660 -20450 4580 -20430
rect 2220 -20510 4580 -20450
rect 30558 -18730 31022 -18560
rect 4060 -20630 4380 -20590
rect 4060 -20770 4100 -20630
rect 4340 -20770 4380 -20630
rect 4060 -20810 4380 -20770
rect 30558 -21304 31020 -18730
rect 30556 -21328 31020 -21304
rect 30556 -21892 31018 -21328
rect 30554 -21920 31018 -21892
rect 30554 -23242 31016 -21920
rect 30552 -23362 31016 -23242
rect 30552 -23516 31014 -23362
rect 30550 -23728 31014 -23516
rect 29280 -23764 31014 -23728
rect 29280 -24096 29318 -23764
rect 29670 -23858 31014 -23764
rect 29670 -24096 31012 -23858
rect 29280 -24130 31012 -24096
<< viali >>
rect 30626 -1356 31016 -1166
rect 30692 -1468 30958 -1432
rect -3640 -3110 -3080 -2930
rect 36326 -4168 36668 -3970
rect 2660 -6690 2740 -6650
rect 3974 -6812 4710 -6768
rect -3610 -9340 -3570 -7000
rect -3530 -9340 -3490 -7000
rect -1370 -9340 -1330 -7000
rect -1280 -9340 -1240 -7000
rect -1200 -9340 -1160 -7000
rect -2820 -11940 -2780 -9600
rect -2780 -11940 -2770 -9600
rect -2730 -11940 -2690 -9600
rect -2650 -11940 -2640 -9600
rect -2640 -11940 -2600 -9600
rect -2280 -11940 -2240 -9600
rect -2200 -11940 -2160 -9600
rect -640 -9340 -600 -7000
rect -560 -9340 -520 -7000
rect -470 -9340 -430 -7000
rect -650 -11940 -610 -9600
rect -610 -11940 -600 -9600
rect -560 -11940 -520 -9600
rect -480 -11940 -470 -9600
rect -470 -11940 -430 -9600
rect 90 -9340 130 -7000
rect 170 -9340 210 -7000
rect 260 -9340 300 -7000
rect 30896 -6852 31016 -6732
rect 2420 -9340 2460 -7000
rect 2500 -9340 2540 -7000
rect 1090 -11940 1130 -9600
rect 1170 -11940 1210 -9600
rect 1530 -11940 1570 -9600
rect 1570 -11940 1580 -9600
rect 1620 -11940 1660 -9600
rect 1700 -11940 1710 -9600
rect 1710 -11940 1750 -9600
rect 36318 -9944 36662 -9812
rect 2608 -12816 2892 -12486
rect 29302 -15148 29806 -14786
rect 30842 -15158 31018 -15018
rect 4100 -15410 4240 -15250
rect 2300 -17790 2660 -15590
rect 4140 -17790 4500 -15590
rect 2300 -20450 2660 -18250
rect 4140 -20430 4500 -18230
rect 4100 -20770 4340 -20630
rect 29318 -24096 29670 -23764
<< metal1 >>
rect 3788 -920 4538 -918
rect 14558 -920 23354 -918
rect 3042 -924 8056 -920
rect 12782 -922 27100 -920
rect 9614 -924 31032 -922
rect 3042 -1166 31032 -924
rect 3042 -1356 30626 -1166
rect 31016 -1356 31032 -1166
rect 3042 -1368 31032 -1356
rect 3042 -1370 18130 -1368
rect 21752 -1370 31032 -1368
rect 3042 -1372 14962 -1370
rect 25684 -1372 28456 -1370
rect 3042 -1374 13644 -1372
rect -3700 -2930 -3020 -2890
rect -3700 -3110 -3640 -2930
rect -3080 -3110 -3020 -2930
rect -3700 -3150 -3020 -3110
rect 3042 -6630 3804 -1374
rect 8296 -1376 13644 -1374
rect 30682 -1432 30968 -1416
rect 30682 -1468 30692 -1432
rect 30958 -1468 30968 -1432
rect 30682 -1828 30968 -1468
rect 4724 -1830 30968 -1828
rect 3962 -2288 30968 -1830
rect 2640 -6650 3800 -6630
rect 2640 -6690 2660 -6650
rect 2740 -6690 3800 -6650
rect 2640 -6710 3800 -6690
rect -3820 -7000 2750 -6970
rect -3820 -9340 -3610 -7000
rect -3570 -9340 -3530 -7000
rect -3490 -9340 -1370 -7000
rect -1330 -9340 -1280 -7000
rect -1240 -9340 -1200 -7000
rect -1160 -9340 -640 -7000
rect -600 -9340 -560 -7000
rect -520 -9340 -470 -7000
rect -430 -9340 90 -7000
rect 130 -9340 170 -7000
rect 210 -9340 260 -7000
rect 300 -9340 2420 -7000
rect 2460 -9340 2500 -7000
rect 2540 -7150 2750 -7000
rect 2540 -9230 2640 -7150
rect 2720 -9230 2750 -7150
rect 2540 -9340 2750 -9230
rect -3820 -9370 2750 -9340
rect -3820 -9590 2750 -9570
rect -3820 -9600 2600 -9590
rect -3820 -11940 -2820 -9600
rect -2770 -11940 -2730 -9600
rect -2690 -11940 -2650 -9600
rect -2600 -11940 -2280 -9600
rect -2240 -11940 -2200 -9600
rect -2160 -11940 -650 -9600
rect -600 -11940 -560 -9600
rect -520 -11940 -480 -9600
rect -430 -11940 1090 -9600
rect 1130 -11940 1170 -9600
rect 1210 -11940 1530 -9600
rect 1580 -11940 1620 -9600
rect 1660 -11940 1700 -9600
rect 1750 -11940 2600 -9600
rect -3820 -11950 2600 -11940
rect 2720 -10660 2750 -9590
rect 2720 -10720 2748 -10660
rect 2720 -11950 2750 -10720
rect -3820 -11970 2750 -11950
rect 1140 -12486 2922 -12458
rect 1140 -12816 2608 -12486
rect 2892 -12816 2922 -12486
rect 1140 -12844 2922 -12816
rect 1140 -27328 1974 -12844
rect 3040 -15090 3800 -6710
rect 3962 -6768 4726 -2288
rect 30784 -3526 31032 -3516
rect 30784 -3780 30796 -3526
rect 31020 -3780 31032 -3526
rect 30784 -3790 31032 -3780
rect 35820 -3790 38180 -1510
rect 36288 -3970 36702 -3936
rect 36288 -4168 36326 -3970
rect 36668 -4168 36702 -3970
rect 3962 -6812 3974 -6768
rect 4710 -6812 4726 -6768
rect 3962 -6824 4726 -6812
rect 4886 -6732 31032 -6606
rect 4886 -6852 30896 -6732
rect 31016 -6852 31032 -6732
rect 4886 -7070 31032 -6852
rect 3866 -7802 5584 -7070
rect 3866 -9508 4630 -7802
rect 3866 -12168 4628 -9508
rect 36288 -9812 36702 -4168
rect 37074 -7088 38180 -3790
rect 36288 -9944 36318 -9812
rect 36662 -9944 36702 -9812
rect 36288 -9966 36702 -9944
rect 29280 -12290 30550 -11886
rect 29442 -14768 29832 -14764
rect 3020 -15210 3800 -15090
rect 29280 -14786 29832 -14768
rect 29280 -15148 29302 -14786
rect 29806 -15148 29832 -14786
rect 29280 -15170 29832 -15148
rect 3020 -15250 4280 -15210
rect 3020 -15410 4100 -15250
rect 4240 -15410 4280 -15250
rect 3020 -15430 4280 -15410
rect 2220 -15590 2760 -15530
rect 2220 -17790 2300 -15590
rect 2660 -17790 2760 -15590
rect 2220 -17850 2760 -17790
rect 2220 -18250 2760 -18170
rect 2220 -20450 2300 -18250
rect 2660 -20450 2760 -18250
rect 2220 -20510 2760 -20450
rect 3020 -20590 3800 -15430
rect 29442 -15512 29832 -15170
rect 30002 -14766 30550 -12290
rect 30002 -14768 30656 -14766
rect 30002 -15018 31032 -14768
rect 30002 -15158 30842 -15018
rect 31018 -15158 31032 -15018
rect 30002 -15170 31032 -15158
rect 30002 -15172 30656 -15170
rect 3020 -20630 4380 -20590
rect 3020 -20770 4100 -20630
rect 4340 -20770 4380 -20630
rect 3020 -20810 4380 -20770
rect 29442 -20850 29834 -15512
rect 29280 -21248 29834 -20850
rect 29280 -21250 29442 -21248
rect 29280 -23764 29712 -23728
rect 29280 -24096 29318 -23764
rect 29670 -24096 29712 -23764
rect 29280 -24130 29712 -24096
rect 1140 -27330 3882 -27328
rect 30642 -27330 31032 -15440
rect 1140 -27790 31032 -27330
rect 1140 -27794 3948 -27790
<< via1 >>
rect -3640 -3110 -3080 -2930
rect 2640 -9230 2720 -7150
rect 2600 -11950 2720 -9590
rect 30796 -3780 31020 -3526
rect 2300 -17790 2660 -15590
rect 2300 -20450 2660 -18250
<< metal2 >>
rect -3700 -2930 -2140 -2890
rect -3700 -3110 -3640 -2930
rect -3080 -3110 -2140 -2930
rect -3700 -15530 -2140 -3110
rect 29012 -3526 31032 -3516
rect 29012 -3780 30796 -3526
rect 31020 -3780 31032 -3526
rect 29012 -3790 31032 -3780
rect 2620 -7150 8260 -7130
rect 2620 -9230 2640 -7150
rect 2720 -8810 8260 -7150
rect 29012 -8810 29280 -3790
rect 2720 -9230 6620 -8810
rect 2620 -9250 6620 -9230
rect 2580 -9590 4060 -9570
rect 2580 -11950 2600 -9590
rect 2720 -11950 4060 -9590
rect 2580 -11970 4060 -11950
rect -3700 -15590 2760 -15530
rect -3700 -17790 2300 -15590
rect 2660 -17790 2760 -15590
rect -3700 -18250 2760 -17790
rect -3700 -20450 2300 -18250
rect 2660 -20450 2760 -18250
rect -3700 -20510 2760 -20450
use bias_gen_resistor  bias_gen_resistor_0
timestamp 1701110497
transform 1 0 -15230 0 1 -12740
box 50 710 11410 12750
use cascode_mirror  cascode_mirror_0
timestamp 1701053371
transform 1 0 38174 0 1 -9726
box -1380 -2940 3780 2640
use ladder_7bit  ladder_7bit_0
timestamp 1701113382
transform 1 0 5320 0 1 -11770
box -1260 -15440 23960 2960
use output_sink  output_sink_0
timestamp 1701111590
transform 1 0 29832 0 1 -13290
box 1200 -4620 6006 12000
<< labels >>
rlabel metal1 -3820 -7710 -3820 -7710 7 VP
port 3 w
rlabel metal1 -3820 -10790 -3820 -10790 7 VN
port 9 w
rlabel locali 2750 -6790 2750 -6790 3 Vcp
port 2 w
rlabel locali -3820 -6670 -3820 -6670 7 Vbp
port 1 w
rlabel locali 2750 -12144 2750 -12144 3 Vcn
port 5 w
<< end >>
