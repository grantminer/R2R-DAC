** sch_path: /home/madvlsi/Documents/R2R-DAC/test_harness_current_mirror.sch
**.subckt test_harness_current_mirror
Vout net1 GND 1
Iref GND net4 100n
XM2 Vbp Vbp VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net3 Vbn GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 Vbn Vbn GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
Vout_i_in net4 Vbn 0
.save i(vout_i_in)
Vout_i_mid Vbp net3 0
.save i(vout_i_mid)
Vout_i_out net2 net1 0
.save i(vout_i_out)
Vdd VDD GND 1.8
**** begin user architecture code


.control
   dc Vout 0 1.8 0.01
   plot i(Vout_i_in) i(Vout_i_mid) i(Vout_i_out)
.endc


.option wnflag=1
.param MC_SWITCH=0.0
.lib ~/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice tt

**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
