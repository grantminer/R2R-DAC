magic
tech sky130A
timestamp 1700691826
<< nwell >>
rect 30 1745 7270 2990
<< nmos >>
rect 450 145 850 1345
rect 2040 145 2440 1345
rect 3270 145 3670 1345
rect 4860 145 5260 1345
<< pmos >>
rect 450 1770 850 2970
rect 2040 1770 2440 2970
rect 3270 1770 3670 2970
rect 4860 1770 5260 2970
rect 6450 1770 6850 2970
<< ndiff >>
rect 50 1285 450 1345
rect 50 205 110 1285
rect 390 205 450 1285
rect 50 145 450 205
rect 850 1285 1250 1345
rect 1640 1285 2040 1345
rect 850 205 910 1285
rect 1190 205 1250 1285
rect 1640 205 1700 1285
rect 1980 205 2040 1285
rect 850 145 1250 205
rect 1640 145 2040 205
rect 2440 1285 2840 1345
rect 2440 205 2500 1285
rect 2780 205 2840 1285
rect 2440 145 2840 205
rect 2870 1285 3270 1345
rect 2870 205 2930 1285
rect 3210 205 3270 1285
rect 2870 145 3270 205
rect 3670 1285 4070 1345
rect 4460 1285 4860 1345
rect 3670 205 3730 1285
rect 4010 205 4070 1285
rect 4460 205 4520 1285
rect 4800 205 4860 1285
rect 3670 145 4070 205
rect 4460 145 4860 205
rect 5260 1285 5660 1345
rect 5260 205 5320 1285
rect 5600 205 5660 1285
rect 5260 145 5660 205
<< pdiff >>
rect 50 2910 450 2970
rect 50 1830 110 2910
rect 390 1830 450 2910
rect 50 1770 450 1830
rect 850 2910 1250 2970
rect 1640 2910 2040 2970
rect 850 1830 910 2910
rect 1190 1830 1250 2910
rect 1640 1830 1700 2910
rect 1980 1830 2040 2910
rect 850 1770 1250 1830
rect 1640 1770 2040 1830
rect 2440 2910 2840 2970
rect 2440 1830 2500 2910
rect 2780 1830 2840 2910
rect 2440 1770 2840 1830
rect 2870 2910 3270 2970
rect 2870 1830 2930 2910
rect 3210 1830 3270 2910
rect 2870 1770 3270 1830
rect 3670 2910 4070 2970
rect 4460 2910 4860 2970
rect 3670 1830 3730 2910
rect 4010 1830 4070 2910
rect 4460 1830 4520 2910
rect 4800 1830 4860 2910
rect 3670 1770 4070 1830
rect 4460 1770 4860 1830
rect 5260 2910 5660 2970
rect 6050 2910 6450 2970
rect 5260 1830 5320 2910
rect 5600 1830 5660 2910
rect 6050 1830 6110 2910
rect 6390 1830 6450 2910
rect 5260 1770 5660 1830
rect 6050 1770 6450 1830
rect 6850 2910 7250 2970
rect 6850 1830 6910 2910
rect 7190 1830 7250 2910
rect 6850 1770 7250 1830
<< ndiffc >>
rect 110 205 390 1285
rect 910 205 1190 1285
rect 1700 205 1980 1285
rect 2500 205 2780 1285
rect 2930 205 3210 1285
rect 3730 205 4010 1285
rect 4520 205 4800 1285
rect 5320 205 5600 1285
<< pdiffc >>
rect 110 1830 390 2910
rect 910 1830 1190 2910
rect 1700 1830 1980 2910
rect 2500 1830 2780 2910
rect 2930 1830 3210 2910
rect 3730 1830 4010 2910
rect 4520 1830 4800 2910
rect 5320 1830 5600 2910
rect 6110 1830 6390 2910
rect 6910 1830 7190 2910
<< psubdiff >>
rect 1250 1285 1640 1345
rect 1250 205 1305 1285
rect 1585 205 1640 1285
rect 1250 145 1640 205
rect 4070 1285 4460 1345
rect 4070 205 4125 1285
rect 4405 205 4460 1285
rect 4070 145 4460 205
<< nsubdiff >>
rect 1250 2910 1640 2970
rect 1250 1830 1305 2910
rect 1585 1830 1640 2910
rect 1250 1770 1640 1830
rect 4070 2910 4460 2970
rect 4070 1830 4125 2910
rect 4405 1830 4460 2910
rect 4070 1770 4460 1830
rect 5660 2910 6050 2970
rect 5660 1830 5715 2910
rect 5995 1830 6050 2910
rect 5660 1770 6050 1830
<< psubdiffcont >>
rect 1305 205 1585 1285
rect 4125 205 4405 1285
<< nsubdiffcont >>
rect 1305 1830 1585 2910
rect 4125 1830 4405 2910
rect 5715 1830 5995 2910
<< poly >>
rect 450 3090 6850 3110
rect 450 3070 3055 3090
rect 3075 3070 6850 3090
rect 450 3060 6850 3070
rect 450 2970 850 3060
rect 2040 2970 2440 3020
rect 3270 2970 3670 3020
rect 4860 2970 5260 3060
rect 6450 2970 6850 3060
rect 450 1720 850 1770
rect 2040 1720 2440 1770
rect 3270 1720 3670 1770
rect 4860 1720 5260 1770
rect 6450 1720 6850 1770
rect 2040 1710 3670 1720
rect 2040 1690 2625 1710
rect 2645 1690 3670 1710
rect 2615 1680 2655 1690
rect 230 1385 2440 1395
rect 5440 1390 5480 1395
rect 230 1365 240 1385
rect 260 1375 2440 1385
rect 260 1365 850 1375
rect 230 1355 850 1365
rect 450 1345 850 1355
rect 2040 1345 2440 1375
rect 3270 1385 5480 1390
rect 3270 1375 5450 1385
rect 3270 1345 3670 1375
rect 4860 1365 5450 1375
rect 5470 1365 5480 1385
rect 4860 1355 5480 1365
rect 4860 1345 5260 1355
rect 450 115 850 145
rect 2040 115 2440 145
rect 3270 115 3670 145
rect 4860 115 5260 145
<< polycont >>
rect 3055 3070 3075 3090
rect 2625 1690 2645 1710
rect 240 1365 260 1385
rect 5450 1365 5470 1385
<< locali >>
rect 3045 3090 3085 3100
rect 3045 3070 3055 3090
rect 3075 3070 3085 3090
rect 230 2940 270 2970
rect 3045 2940 3085 3070
rect 5440 2940 5480 2970
rect 7030 2940 7070 2970
rect 80 2910 420 2940
rect 80 1830 110 2910
rect 390 1830 420 2910
rect 80 1800 420 1830
rect 880 2910 2010 2940
rect 880 1830 910 2910
rect 1190 1830 1305 2910
rect 1585 1830 1700 2910
rect 1980 1830 2010 2910
rect 880 1805 2010 1830
rect 1300 1800 2010 1805
rect 2470 2910 2810 2940
rect 2470 1830 2500 2910
rect 2780 1830 2810 2910
rect 2470 1710 2810 1830
rect 2470 1690 2625 1710
rect 2645 1690 2810 1710
rect 230 1385 270 1395
rect 230 1365 240 1385
rect 260 1365 270 1385
rect 230 1315 270 1365
rect 80 1285 420 1315
rect 80 205 110 1285
rect 390 205 420 1285
rect 80 175 420 205
rect 880 1285 1220 1315
rect 880 205 910 1285
rect 1190 205 1220 1285
rect 880 -105 1220 205
rect 1275 1285 2010 1315
rect 1275 205 1305 1285
rect 1585 205 1700 1285
rect 1980 205 2010 1285
rect 1275 175 2010 205
rect 2470 1285 2810 1690
rect 2470 205 2500 1285
rect 2780 205 2810 1285
rect 2470 175 2810 205
rect 2900 2910 3240 2940
rect 2900 1830 2930 2910
rect 3210 1830 3240 2910
rect 2900 1285 3240 1830
rect 3700 2910 4830 2940
rect 3700 1830 3730 2910
rect 4010 1830 4125 2910
rect 4405 1830 4520 2910
rect 4800 1830 4830 2910
rect 3700 1800 4830 1830
rect 5290 2910 5630 2940
rect 5290 1830 5320 2910
rect 5600 1830 5630 2910
rect 5290 1800 5630 1830
rect 5660 2910 6420 2940
rect 5660 1830 5715 2910
rect 5995 1830 6110 2910
rect 6390 1830 6420 2910
rect 5660 1800 6420 1830
rect 6880 2910 7220 2940
rect 6880 1830 6910 2910
rect 7190 1830 7220 2910
rect 6880 1800 7220 1830
rect 5440 1385 5480 1395
rect 5440 1365 5450 1385
rect 5470 1365 5480 1385
rect 5440 1315 5480 1365
rect 2900 205 2930 1285
rect 3210 205 3240 1285
rect 2900 175 3240 205
rect 3700 1285 4830 1315
rect 3700 205 3730 1285
rect 4010 205 4125 1285
rect 4405 205 4520 1285
rect 4800 205 4830 1285
rect 3700 175 4830 205
rect 5290 1285 5630 1315
rect 5290 205 5320 1285
rect 5600 205 5630 1285
rect 5290 175 5630 205
<< labels >>
flabel space 855 -380 1150 0 0 FreeSans 800 0 0 0 R
flabel pmos 475 1795 770 2175 0 FreeSans 800 0 0 0 VG
<< end >>
