magic
tech sky130A
timestamp 1701150901
<< nwell >>
rect 630 -20 2300 1220
rect 4010 -20 5680 1220
rect 7390 -20 9060 1220
rect 10770 -20 11700 1220
rect 630 -7460 2300 -6220
rect 4010 -7460 5680 -6220
rect 7390 -7460 9060 -6220
rect 10770 -7460 11700 -6220
<< nmos >>
rect 0 0 400 1200
rect 2530 0 2930 1200
rect 3380 0 3780 1200
rect 5910 0 6310 1200
rect 6760 0 7160 1200
rect 9290 0 9690 1200
rect 10140 0 10540 1200
rect 0 -1480 400 -280
rect 840 -1480 1240 -280
rect 1690 -1480 2090 -280
rect 2530 -1480 2930 -280
rect 3380 -1480 3780 -280
rect 4220 -1480 4620 -280
rect 5070 -1480 5470 -280
rect 5910 -1480 6310 -280
rect 6760 -1480 7160 -280
rect 7600 -1480 8000 -280
rect 8450 -1480 8850 -280
rect 9290 -1480 9690 -280
rect 10140 -1480 10540 -280
rect 10980 -1480 11380 -280
rect 0 -3060 400 -1860
rect 840 -3060 1240 -1860
rect 1690 -3060 2090 -1860
rect 2530 -3060 2930 -1860
rect 3380 -3060 3780 -1860
rect 4220 -3060 4620 -1860
rect 5070 -3060 5470 -1860
rect 5910 -3060 6310 -1860
rect 6760 -3060 7160 -1860
rect 7600 -3060 8000 -1860
rect 8450 -3060 8850 -1860
rect 9290 -3060 9690 -1860
rect 10140 -3060 10540 -1860
rect 10980 -3060 11380 -1860
rect 11420 -3060 11820 -1860
rect 0 -4380 400 -3180
rect 840 -4380 1240 -3180
rect 1690 -4380 2090 -3180
rect 2530 -4380 2930 -3180
rect 3380 -4380 3780 -3180
rect 4220 -4380 4620 -3180
rect 5070 -4380 5470 -3180
rect 5910 -4380 6310 -3180
rect 6760 -4380 7160 -3180
rect 7600 -4380 8000 -3180
rect 8450 -4380 8850 -3180
rect 9290 -4380 9690 -3180
rect 10140 -4380 10540 -3180
rect 10980 -4380 11380 -3180
rect 11420 -4380 11820 -3180
rect 0 -5960 400 -4760
rect 840 -5960 1240 -4760
rect 1690 -5960 2090 -4760
rect 2530 -5960 2930 -4760
rect 3380 -5960 3780 -4760
rect 4220 -5960 4620 -4760
rect 5070 -5960 5470 -4760
rect 5910 -5960 6310 -4760
rect 6760 -5960 7160 -4760
rect 7600 -5960 8000 -4760
rect 8450 -5960 8850 -4760
rect 9290 -5960 9690 -4760
rect 10140 -5960 10540 -4760
rect 10980 -5960 11380 -4760
rect 0 -7440 400 -6240
rect 2530 -7440 2930 -6240
rect 3380 -7440 3780 -6240
rect 5910 -7440 6310 -6240
rect 6760 -7440 7160 -6240
rect 9290 -7440 9690 -6240
rect 10140 -7440 10540 -6240
<< pmos >>
rect 840 0 1240 1200
rect 1690 0 2090 1200
rect 4220 0 4620 1200
rect 5070 0 5470 1200
rect 7600 0 8000 1200
rect 8450 0 8850 1200
rect 10980 0 11380 1200
rect 840 -7440 1240 -6240
rect 1690 -7440 2090 -6240
rect 4220 -7440 4620 -6240
rect 5070 -7440 5470 -6240
rect 7600 -7440 8000 -6240
rect 8450 -7440 8850 -6240
rect 10980 -7440 11380 -6240
<< ndiff >>
rect -160 1140 0 1200
rect -160 60 -130 1140
rect -60 60 0 1140
rect -160 0 0 60
rect 400 1130 590 1200
rect 400 60 460 1130
rect 530 60 590 1130
rect 400 0 590 60
rect 2340 1130 2530 1200
rect 2340 60 2400 1130
rect 2470 60 2530 1130
rect 2340 0 2530 60
rect 2930 1140 3090 1200
rect 3220 1140 3380 1200
rect 2930 60 2990 1140
rect 3060 60 3090 1140
rect 3220 60 3250 1140
rect 3320 60 3380 1140
rect 2930 0 3090 60
rect 3220 0 3380 60
rect 3780 1130 3970 1200
rect 3780 60 3840 1130
rect 3910 60 3970 1130
rect 3780 0 3970 60
rect 5720 1130 5910 1200
rect 5720 60 5780 1130
rect 5850 60 5910 1130
rect 5720 0 5910 60
rect 6310 1140 6470 1200
rect 6600 1140 6760 1200
rect 6310 60 6370 1140
rect 6440 60 6470 1140
rect 6600 60 6630 1140
rect 6700 60 6760 1140
rect 6310 0 6470 60
rect 6600 0 6760 60
rect 7160 1130 7350 1200
rect 7160 60 7220 1130
rect 7290 60 7350 1130
rect 7160 0 7350 60
rect 9100 1130 9290 1200
rect 9100 60 9160 1130
rect 9230 60 9290 1130
rect 9100 0 9290 60
rect 9690 1140 9850 1200
rect 9980 1140 10140 1200
rect 9690 60 9750 1140
rect 9820 60 9850 1140
rect 9980 60 10010 1140
rect 10080 60 10140 1140
rect 9690 0 9850 60
rect 9980 0 10140 60
rect 10540 1130 10730 1200
rect 10540 60 10600 1130
rect 10670 60 10730 1130
rect 10540 0 10730 60
rect -160 -320 0 -280
rect -160 -1440 -120 -320
rect -40 -1440 0 -320
rect -160 -1480 0 -1440
rect 400 -340 840 -280
rect 400 -1420 460 -340
rect 780 -1420 840 -340
rect 400 -1480 840 -1420
rect 1240 -320 1400 -280
rect 1240 -1440 1280 -320
rect 1360 -1440 1400 -320
rect 1240 -1480 1400 -1440
rect 1530 -320 1690 -280
rect 1530 -1440 1570 -320
rect 1650 -1440 1690 -320
rect 1530 -1480 1690 -1440
rect 2090 -340 2530 -280
rect 2090 -1420 2150 -340
rect 2470 -1420 2530 -340
rect 2090 -1480 2530 -1420
rect 2930 -320 3090 -280
rect 2930 -1440 2970 -320
rect 3050 -1440 3090 -320
rect 2930 -1480 3090 -1440
rect 3220 -320 3380 -280
rect 3220 -1440 3260 -320
rect 3340 -1440 3380 -320
rect 3220 -1480 3380 -1440
rect 3780 -340 4220 -280
rect 3780 -1420 3840 -340
rect 4160 -1420 4220 -340
rect 3780 -1480 4220 -1420
rect 4620 -320 4780 -280
rect 4620 -1440 4660 -320
rect 4740 -1440 4780 -320
rect 4620 -1480 4780 -1440
rect 4910 -320 5070 -280
rect 4910 -1440 4950 -320
rect 5030 -1440 5070 -320
rect 4910 -1480 5070 -1440
rect 5470 -340 5910 -280
rect 5470 -1420 5530 -340
rect 5850 -1420 5910 -340
rect 5470 -1480 5910 -1420
rect 6310 -320 6470 -280
rect 6310 -1440 6350 -320
rect 6430 -1440 6470 -320
rect 6310 -1480 6470 -1440
rect 6600 -320 6760 -280
rect 6600 -1440 6640 -320
rect 6720 -1440 6760 -320
rect 6600 -1480 6760 -1440
rect 7160 -340 7600 -280
rect 7160 -1420 7220 -340
rect 7540 -1420 7600 -340
rect 7160 -1480 7600 -1420
rect 8000 -320 8160 -280
rect 8000 -1440 8040 -320
rect 8120 -1440 8160 -320
rect 8000 -1480 8160 -1440
rect 8290 -320 8450 -280
rect 8290 -1440 8330 -320
rect 8410 -1440 8450 -320
rect 8290 -1480 8450 -1440
rect 8850 -340 9290 -280
rect 8850 -1420 8910 -340
rect 9230 -1420 9290 -340
rect 8850 -1480 9290 -1420
rect 9690 -320 9850 -280
rect 9690 -1440 9730 -320
rect 9810 -1440 9850 -320
rect 9690 -1480 9850 -1440
rect 9980 -320 10140 -280
rect 9980 -1440 10020 -320
rect 10100 -1440 10140 -320
rect 9980 -1480 10140 -1440
rect 10540 -340 10980 -280
rect 10540 -1420 10600 -340
rect 10920 -1420 10980 -340
rect 10540 -1480 10980 -1420
rect 11380 -320 11540 -280
rect 11380 -1440 11420 -320
rect 11500 -1440 11540 -320
rect 11380 -1480 11540 -1440
rect -160 -1900 0 -1860
rect -160 -3020 -120 -1900
rect -40 -3020 0 -1900
rect -160 -3060 0 -3020
rect 400 -1910 840 -1860
rect 400 -3010 460 -1910
rect 780 -3010 840 -1910
rect 400 -3060 840 -3010
rect 1240 -1900 1400 -1860
rect 1240 -3020 1280 -1900
rect 1360 -3020 1400 -1900
rect 1240 -3060 1400 -3020
rect 1530 -1900 1690 -1860
rect 1530 -3020 1570 -1900
rect 1650 -3020 1690 -1900
rect 1530 -3060 1690 -3020
rect 2090 -1910 2530 -1860
rect 2090 -3010 2150 -1910
rect 2470 -3010 2530 -1910
rect 2090 -3060 2530 -3010
rect 2930 -1900 3090 -1860
rect 2930 -3020 2970 -1900
rect 3050 -3020 3090 -1900
rect 2930 -3060 3090 -3020
rect 3220 -1900 3380 -1860
rect 3220 -3020 3260 -1900
rect 3340 -3020 3380 -1900
rect 3220 -3060 3380 -3020
rect 3780 -1910 4220 -1860
rect 3780 -3010 3840 -1910
rect 4160 -3010 4220 -1910
rect 3780 -3060 4220 -3010
rect 4620 -1900 4780 -1860
rect 4620 -3020 4660 -1900
rect 4740 -3020 4780 -1900
rect 4620 -3060 4780 -3020
rect 4910 -1900 5070 -1860
rect 4910 -3020 4950 -1900
rect 5030 -3020 5070 -1900
rect 4910 -3060 5070 -3020
rect 5470 -1910 5910 -1860
rect 5470 -3010 5530 -1910
rect 5850 -3010 5910 -1910
rect 5470 -3060 5910 -3010
rect 6310 -1900 6470 -1860
rect 6310 -3020 6350 -1900
rect 6430 -3020 6470 -1900
rect 6310 -3060 6470 -3020
rect 6600 -1900 6760 -1860
rect 6600 -3020 6640 -1900
rect 6720 -3020 6760 -1900
rect 6600 -3060 6760 -3020
rect 7160 -1910 7600 -1860
rect 7160 -3010 7220 -1910
rect 7540 -3010 7600 -1910
rect 7160 -3060 7600 -3010
rect 8000 -1900 8160 -1860
rect 8000 -3020 8040 -1900
rect 8120 -3020 8160 -1900
rect 8000 -3060 8160 -3020
rect 8290 -1900 8450 -1860
rect 8290 -3020 8330 -1900
rect 8410 -3020 8450 -1900
rect 8290 -3060 8450 -3020
rect 8850 -1910 9290 -1860
rect 8850 -3010 8910 -1910
rect 9230 -3010 9290 -1910
rect 8850 -3060 9290 -3010
rect 9690 -1900 9850 -1860
rect 9690 -3020 9730 -1900
rect 9810 -3020 9850 -1900
rect 9690 -3060 9850 -3020
rect 9980 -1900 10140 -1860
rect 9980 -3020 10020 -1900
rect 10100 -3020 10140 -1900
rect 9980 -3060 10140 -3020
rect 10540 -1910 10980 -1860
rect 10540 -3010 10600 -1910
rect 10920 -3010 10980 -1910
rect 10540 -3060 10980 -3010
rect 11380 -3060 11420 -1860
rect 11820 -1900 11980 -1860
rect 11820 -3020 11860 -1900
rect 11940 -3020 11980 -1900
rect 11820 -3060 11980 -3020
rect -160 -3220 0 -3180
rect -160 -4340 -120 -3220
rect -40 -4340 0 -3220
rect -160 -4380 0 -4340
rect 400 -3230 840 -3180
rect 400 -4330 460 -3230
rect 780 -4330 840 -3230
rect 400 -4380 840 -4330
rect 1240 -3220 1400 -3180
rect 1240 -4340 1280 -3220
rect 1360 -4340 1400 -3220
rect 1240 -4380 1400 -4340
rect 1530 -3220 1690 -3180
rect 1530 -4340 1570 -3220
rect 1650 -4340 1690 -3220
rect 1530 -4380 1690 -4340
rect 2090 -3230 2530 -3180
rect 2090 -4330 2150 -3230
rect 2470 -4330 2530 -3230
rect 2090 -4380 2530 -4330
rect 2930 -3220 3090 -3180
rect 2930 -4340 2970 -3220
rect 3050 -4340 3090 -3220
rect 2930 -4380 3090 -4340
rect 3220 -3220 3380 -3180
rect 3220 -4340 3260 -3220
rect 3340 -4340 3380 -3220
rect 3220 -4380 3380 -4340
rect 3780 -3230 4220 -3180
rect 3780 -4330 3840 -3230
rect 4160 -4330 4220 -3230
rect 3780 -4380 4220 -4330
rect 4620 -3220 4780 -3180
rect 4620 -4340 4660 -3220
rect 4740 -4340 4780 -3220
rect 4620 -4380 4780 -4340
rect 4910 -3220 5070 -3180
rect 4910 -4340 4950 -3220
rect 5030 -4340 5070 -3220
rect 4910 -4380 5070 -4340
rect 5470 -3230 5910 -3180
rect 5470 -4330 5530 -3230
rect 5850 -4330 5910 -3230
rect 5470 -4380 5910 -4330
rect 6310 -3220 6470 -3180
rect 6310 -4340 6350 -3220
rect 6430 -4340 6470 -3220
rect 6310 -4380 6470 -4340
rect 6600 -3220 6760 -3180
rect 6600 -4340 6640 -3220
rect 6720 -4340 6760 -3220
rect 6600 -4380 6760 -4340
rect 7160 -3230 7600 -3180
rect 7160 -4330 7220 -3230
rect 7540 -4330 7600 -3230
rect 7160 -4380 7600 -4330
rect 8000 -3220 8160 -3180
rect 8000 -4340 8040 -3220
rect 8120 -4340 8160 -3220
rect 8000 -4380 8160 -4340
rect 8290 -3220 8450 -3180
rect 8290 -4340 8330 -3220
rect 8410 -4340 8450 -3220
rect 8290 -4380 8450 -4340
rect 8850 -3230 9290 -3180
rect 8850 -4330 8910 -3230
rect 9230 -4330 9290 -3230
rect 8850 -4380 9290 -4330
rect 9690 -3220 9850 -3180
rect 9690 -4340 9730 -3220
rect 9810 -4340 9850 -3220
rect 9690 -4380 9850 -4340
rect 9980 -3220 10140 -3180
rect 9980 -4340 10020 -3220
rect 10100 -4340 10140 -3220
rect 9980 -4380 10140 -4340
rect 10540 -3230 10980 -3180
rect 10540 -4330 10600 -3230
rect 10920 -4330 10980 -3230
rect 10540 -4380 10980 -4330
rect 11380 -4380 11420 -3180
rect 11820 -3220 11980 -3180
rect 11820 -4340 11860 -3220
rect 11940 -4340 11980 -3220
rect 11820 -4380 11980 -4340
rect -160 -4800 0 -4760
rect -160 -5920 -120 -4800
rect -40 -5920 0 -4800
rect -160 -5960 0 -5920
rect 400 -4820 840 -4760
rect 400 -5900 460 -4820
rect 780 -5900 840 -4820
rect 400 -5960 840 -5900
rect 1240 -4800 1400 -4760
rect 1240 -5920 1280 -4800
rect 1360 -5920 1400 -4800
rect 1240 -5960 1400 -5920
rect 1530 -4800 1690 -4760
rect 1530 -5920 1570 -4800
rect 1650 -5920 1690 -4800
rect 1530 -5960 1690 -5920
rect 2090 -4820 2530 -4760
rect 2090 -5900 2150 -4820
rect 2470 -5900 2530 -4820
rect 2090 -5960 2530 -5900
rect 2930 -4800 3090 -4760
rect 2930 -5920 2970 -4800
rect 3050 -5920 3090 -4800
rect 2930 -5960 3090 -5920
rect 3220 -4800 3380 -4760
rect 3220 -5920 3260 -4800
rect 3340 -5920 3380 -4800
rect 3220 -5960 3380 -5920
rect 3780 -4820 4220 -4760
rect 3780 -5900 3840 -4820
rect 4160 -5900 4220 -4820
rect 3780 -5960 4220 -5900
rect 4620 -4800 4780 -4760
rect 4620 -5920 4660 -4800
rect 4740 -5920 4780 -4800
rect 4620 -5960 4780 -5920
rect 4910 -4800 5070 -4760
rect 4910 -5920 4950 -4800
rect 5030 -5920 5070 -4800
rect 4910 -5960 5070 -5920
rect 5470 -4820 5910 -4760
rect 5470 -5900 5530 -4820
rect 5850 -5900 5910 -4820
rect 5470 -5960 5910 -5900
rect 6310 -4800 6470 -4760
rect 6310 -5920 6350 -4800
rect 6430 -5920 6470 -4800
rect 6310 -5960 6470 -5920
rect 6600 -4800 6760 -4760
rect 6600 -5920 6640 -4800
rect 6720 -5920 6760 -4800
rect 6600 -5960 6760 -5920
rect 7160 -4820 7600 -4760
rect 7160 -5900 7220 -4820
rect 7540 -5900 7600 -4820
rect 7160 -5960 7600 -5900
rect 8000 -4800 8160 -4760
rect 8000 -5920 8040 -4800
rect 8120 -5920 8160 -4800
rect 8000 -5960 8160 -5920
rect 8290 -4800 8450 -4760
rect 8290 -5920 8330 -4800
rect 8410 -5920 8450 -4800
rect 8290 -5960 8450 -5920
rect 8850 -4820 9290 -4760
rect 8850 -5900 8910 -4820
rect 9230 -5900 9290 -4820
rect 8850 -5960 9290 -5900
rect 9690 -4800 9850 -4760
rect 9690 -5920 9730 -4800
rect 9810 -5920 9850 -4800
rect 9690 -5960 9850 -5920
rect 9980 -4800 10140 -4760
rect 9980 -5920 10020 -4800
rect 10100 -5920 10140 -4800
rect 9980 -5960 10140 -5920
rect 10540 -4820 10980 -4760
rect 10540 -5900 10600 -4820
rect 10920 -5900 10980 -4820
rect 10540 -5960 10980 -5900
rect 11380 -4800 11540 -4760
rect 11380 -5920 11420 -4800
rect 11500 -5920 11540 -4800
rect 11380 -5960 11540 -5920
rect -160 -6300 0 -6240
rect -160 -7380 -130 -6300
rect -60 -7380 0 -6300
rect -160 -7440 0 -7380
rect 400 -6300 590 -6240
rect 400 -7370 460 -6300
rect 530 -7370 590 -6300
rect 400 -7440 590 -7370
rect 2340 -6300 2530 -6240
rect 2340 -7370 2400 -6300
rect 2470 -7370 2530 -6300
rect 2340 -7440 2530 -7370
rect 2930 -6300 3090 -6240
rect 3220 -6300 3380 -6240
rect 2930 -7380 2990 -6300
rect 3060 -7380 3090 -6300
rect 3220 -7380 3250 -6300
rect 3320 -7380 3380 -6300
rect 2930 -7440 3090 -7380
rect 3220 -7440 3380 -7380
rect 3780 -6300 3970 -6240
rect 3780 -7370 3840 -6300
rect 3910 -7370 3970 -6300
rect 3780 -7440 3970 -7370
rect 5720 -6300 5910 -6240
rect 5720 -7370 5780 -6300
rect 5850 -7370 5910 -6300
rect 5720 -7440 5910 -7370
rect 6310 -6300 6470 -6240
rect 6600 -6300 6760 -6240
rect 6310 -7380 6370 -6300
rect 6440 -7380 6470 -6300
rect 6600 -7380 6630 -6300
rect 6700 -7380 6760 -6300
rect 6310 -7440 6470 -7380
rect 6600 -7440 6760 -7380
rect 7160 -6300 7350 -6240
rect 7160 -7370 7220 -6300
rect 7290 -7370 7350 -6300
rect 7160 -7440 7350 -7370
rect 9100 -6300 9290 -6240
rect 9100 -7370 9160 -6300
rect 9230 -7370 9290 -6300
rect 9100 -7440 9290 -7370
rect 9690 -6300 9850 -6240
rect 9980 -6300 10140 -6240
rect 9690 -7380 9750 -6300
rect 9820 -7380 9850 -6300
rect 9980 -7380 10010 -6300
rect 10080 -7380 10140 -6300
rect 9690 -7440 9850 -7380
rect 9980 -7440 10140 -7380
rect 10540 -6300 10730 -6240
rect 10540 -7370 10600 -6300
rect 10670 -7370 10730 -6300
rect 10540 -7440 10730 -7370
<< pdiff >>
rect 650 1130 840 1200
rect 650 60 710 1130
rect 780 60 840 1130
rect 650 0 840 60
rect 1240 1140 1400 1200
rect 1530 1140 1690 1200
rect 1240 60 1300 1140
rect 1370 60 1400 1140
rect 1530 60 1560 1140
rect 1630 60 1690 1140
rect 1240 0 1400 60
rect 1530 0 1690 60
rect 2090 1130 2280 1200
rect 2090 60 2150 1130
rect 2220 60 2280 1130
rect 2090 0 2280 60
rect 4030 1130 4220 1200
rect 4030 60 4090 1130
rect 4160 60 4220 1130
rect 4030 0 4220 60
rect 4620 1140 4780 1200
rect 4910 1140 5070 1200
rect 4620 60 4680 1140
rect 4750 60 4780 1140
rect 4910 60 4940 1140
rect 5010 60 5070 1140
rect 4620 0 4780 60
rect 4910 0 5070 60
rect 5470 1130 5660 1200
rect 5470 60 5530 1130
rect 5600 60 5660 1130
rect 5470 0 5660 60
rect 7410 1130 7600 1200
rect 7410 60 7470 1130
rect 7540 60 7600 1130
rect 7410 0 7600 60
rect 8000 1140 8160 1200
rect 8290 1140 8450 1200
rect 8000 60 8060 1140
rect 8130 60 8160 1140
rect 8290 60 8320 1140
rect 8390 60 8450 1140
rect 8000 0 8160 60
rect 8290 0 8450 60
rect 8850 1130 9040 1200
rect 8850 60 8910 1130
rect 8980 60 9040 1130
rect 8850 0 9040 60
rect 10790 1130 10980 1200
rect 10790 60 10850 1130
rect 10920 60 10980 1130
rect 10790 0 10980 60
rect 11380 1140 11540 1200
rect 11380 60 11440 1140
rect 11510 60 11540 1140
rect 11380 0 11540 60
rect 650 -6300 840 -6240
rect 650 -7370 710 -6300
rect 780 -7370 840 -6300
rect 650 -7440 840 -7370
rect 1240 -6300 1400 -6240
rect 1530 -6300 1690 -6240
rect 1240 -7380 1300 -6300
rect 1370 -7380 1400 -6300
rect 1530 -7380 1560 -6300
rect 1630 -7380 1690 -6300
rect 1240 -7440 1400 -7380
rect 1530 -7440 1690 -7380
rect 2090 -6300 2280 -6240
rect 2090 -7370 2150 -6300
rect 2220 -7370 2280 -6300
rect 2090 -7440 2280 -7370
rect 4030 -6300 4220 -6240
rect 4030 -7370 4090 -6300
rect 4160 -7370 4220 -6300
rect 4030 -7440 4220 -7370
rect 4620 -6300 4780 -6240
rect 4910 -6300 5070 -6240
rect 4620 -7380 4680 -6300
rect 4750 -7380 4780 -6300
rect 4910 -7380 4940 -6300
rect 5010 -7380 5070 -6300
rect 4620 -7440 4780 -7380
rect 4910 -7440 5070 -7380
rect 5470 -6300 5660 -6240
rect 5470 -7370 5530 -6300
rect 5600 -7370 5660 -6300
rect 5470 -7440 5660 -7370
rect 7410 -6300 7600 -6240
rect 7410 -7370 7470 -6300
rect 7540 -7370 7600 -6300
rect 7410 -7440 7600 -7370
rect 8000 -6300 8160 -6240
rect 8290 -6300 8450 -6240
rect 8000 -7380 8060 -6300
rect 8130 -7380 8160 -6300
rect 8290 -7380 8320 -6300
rect 8390 -7380 8450 -6300
rect 8000 -7440 8160 -7380
rect 8290 -7440 8450 -7380
rect 8850 -6300 9040 -6240
rect 8850 -7370 8910 -6300
rect 8980 -7370 9040 -6300
rect 8850 -7440 9040 -7370
rect 10790 -6300 10980 -6240
rect 10790 -7370 10850 -6300
rect 10920 -7370 10980 -6300
rect 10790 -7440 10980 -7370
rect 11380 -6300 11540 -6240
rect 11380 -7380 11440 -6300
rect 11510 -7380 11540 -6300
rect 11380 -7440 11540 -7380
<< ndiffc >>
rect -130 60 -60 1140
rect 460 60 530 1130
rect 2400 60 2470 1130
rect 2990 60 3060 1140
rect 3250 60 3320 1140
rect 3840 60 3910 1130
rect 5780 60 5850 1130
rect 6370 60 6440 1140
rect 6630 60 6700 1140
rect 7220 60 7290 1130
rect 9160 60 9230 1130
rect 9750 60 9820 1140
rect 10010 60 10080 1140
rect 10600 60 10670 1130
rect -120 -1440 -40 -320
rect 460 -1420 780 -340
rect 1280 -1440 1360 -320
rect 1570 -1440 1650 -320
rect 2150 -1420 2470 -340
rect 2970 -1440 3050 -320
rect 3260 -1440 3340 -320
rect 3840 -1420 4160 -340
rect 4660 -1440 4740 -320
rect 4950 -1440 5030 -320
rect 5530 -1420 5850 -340
rect 6350 -1440 6430 -320
rect 6640 -1440 6720 -320
rect 7220 -1420 7540 -340
rect 8040 -1440 8120 -320
rect 8330 -1440 8410 -320
rect 8910 -1420 9230 -340
rect 9730 -1440 9810 -320
rect 10020 -1440 10100 -320
rect 10600 -1420 10920 -340
rect 11420 -1440 11500 -320
rect -120 -3020 -40 -1900
rect 460 -3010 780 -1910
rect 1280 -3020 1360 -1900
rect 1570 -3020 1650 -1900
rect 2150 -3010 2470 -1910
rect 2970 -3020 3050 -1900
rect 3260 -3020 3340 -1900
rect 3840 -3010 4160 -1910
rect 4660 -3020 4740 -1900
rect 4950 -3020 5030 -1900
rect 5530 -3010 5850 -1910
rect 6350 -3020 6430 -1900
rect 6640 -3020 6720 -1900
rect 7220 -3010 7540 -1910
rect 8040 -3020 8120 -1900
rect 8330 -3020 8410 -1900
rect 8910 -3010 9230 -1910
rect 9730 -3020 9810 -1900
rect 10020 -3020 10100 -1900
rect 10600 -3010 10920 -1910
rect 11860 -3020 11940 -1900
rect -120 -4340 -40 -3220
rect 460 -4330 780 -3230
rect 1280 -4340 1360 -3220
rect 1570 -4340 1650 -3220
rect 2150 -4330 2470 -3230
rect 2970 -4340 3050 -3220
rect 3260 -4340 3340 -3220
rect 3840 -4330 4160 -3230
rect 4660 -4340 4740 -3220
rect 4950 -4340 5030 -3220
rect 5530 -4330 5850 -3230
rect 6350 -4340 6430 -3220
rect 6640 -4340 6720 -3220
rect 7220 -4330 7540 -3230
rect 8040 -4340 8120 -3220
rect 8330 -4340 8410 -3220
rect 8910 -4330 9230 -3230
rect 9730 -4340 9810 -3220
rect 10020 -4340 10100 -3220
rect 10600 -4330 10920 -3230
rect 11860 -4340 11940 -3220
rect -120 -5920 -40 -4800
rect 460 -5900 780 -4820
rect 1280 -5920 1360 -4800
rect 1570 -5920 1650 -4800
rect 2150 -5900 2470 -4820
rect 2970 -5920 3050 -4800
rect 3260 -5920 3340 -4800
rect 3840 -5900 4160 -4820
rect 4660 -5920 4740 -4800
rect 4950 -5920 5030 -4800
rect 5530 -5900 5850 -4820
rect 6350 -5920 6430 -4800
rect 6640 -5920 6720 -4800
rect 7220 -5900 7540 -4820
rect 8040 -5920 8120 -4800
rect 8330 -5920 8410 -4800
rect 8910 -5900 9230 -4820
rect 9730 -5920 9810 -4800
rect 10020 -5920 10100 -4800
rect 10600 -5900 10920 -4820
rect 11420 -5920 11500 -4800
rect -130 -7380 -60 -6300
rect 460 -7370 530 -6300
rect 2400 -7370 2470 -6300
rect 2990 -7380 3060 -6300
rect 3250 -7380 3320 -6300
rect 3840 -7370 3910 -6300
rect 5780 -7370 5850 -6300
rect 6370 -7380 6440 -6300
rect 6630 -7380 6700 -6300
rect 7220 -7370 7290 -6300
rect 9160 -7370 9230 -6300
rect 9750 -7380 9820 -6300
rect 10010 -7380 10080 -6300
rect 10600 -7370 10670 -6300
<< pdiffc >>
rect 710 60 780 1130
rect 1300 60 1370 1140
rect 1560 60 1630 1140
rect 2150 60 2220 1130
rect 4090 60 4160 1130
rect 4680 60 4750 1140
rect 4940 60 5010 1140
rect 5530 60 5600 1130
rect 7470 60 7540 1130
rect 8060 60 8130 1140
rect 8320 60 8390 1140
rect 8910 60 8980 1130
rect 10850 60 10920 1130
rect 11440 60 11510 1140
rect 710 -7370 780 -6300
rect 1300 -7380 1370 -6300
rect 1560 -7380 1630 -6300
rect 2150 -7370 2220 -6300
rect 4090 -7370 4160 -6300
rect 4680 -7380 4750 -6300
rect 4940 -7380 5010 -6300
rect 5530 -7370 5600 -6300
rect 7470 -7370 7540 -6300
rect 8060 -7380 8130 -6300
rect 8320 -7380 8390 -6300
rect 8910 -7370 8980 -6300
rect 10850 -7370 10920 -6300
rect 11440 -7380 11510 -6300
<< psubdiff >>
rect -330 1140 -160 1200
rect -330 60 -290 1140
rect -190 60 -160 1140
rect -330 0 -160 60
rect 3090 1140 3220 1200
rect 3090 60 3120 1140
rect 3190 60 3220 1140
rect 3090 0 3220 60
rect 6470 1140 6600 1200
rect 6470 60 6500 1140
rect 6570 60 6600 1140
rect 6470 0 6600 60
rect 9850 1140 9980 1200
rect 9850 60 9880 1140
rect 9950 60 9980 1140
rect 9850 0 9980 60
rect -330 -6300 -160 -6240
rect -330 -7380 -290 -6300
rect -190 -7380 -160 -6300
rect -330 -7440 -160 -7380
rect 3090 -6300 3220 -6240
rect 3090 -7380 3120 -6300
rect 3190 -7380 3220 -6300
rect 3090 -7440 3220 -7380
rect 6470 -6300 6600 -6240
rect 6470 -7380 6500 -6300
rect 6570 -7380 6600 -6300
rect 6470 -7440 6600 -7380
rect 9850 -6300 9980 -6240
rect 9850 -7380 9880 -6300
rect 9950 -7380 9980 -6300
rect 9850 -7440 9980 -7380
<< nsubdiff >>
rect 1400 1140 1530 1200
rect 1400 60 1430 1140
rect 1500 60 1530 1140
rect 1400 0 1530 60
rect 4780 1140 4910 1200
rect 4780 60 4810 1140
rect 4880 60 4910 1140
rect 4780 0 4910 60
rect 8160 1140 8290 1200
rect 8160 60 8190 1140
rect 8260 60 8290 1140
rect 8160 0 8290 60
rect 11540 1140 11680 1200
rect 11540 60 11570 1140
rect 11640 60 11680 1140
rect 11540 0 11680 60
rect 1400 -6300 1530 -6240
rect 1400 -7380 1430 -6300
rect 1500 -7380 1530 -6300
rect 1400 -7440 1530 -7380
rect 4780 -6300 4910 -6240
rect 4780 -7380 4810 -6300
rect 4880 -7380 4910 -6300
rect 4780 -7440 4910 -7380
rect 8160 -6300 8290 -6240
rect 8160 -7380 8190 -6300
rect 8260 -7380 8290 -6300
rect 8160 -7440 8290 -7380
rect 11540 -6300 11680 -6240
rect 11540 -7380 11570 -6300
rect 11640 -7380 11680 -6300
rect 11540 -7440 11680 -7380
<< psubdiffcont >>
rect -290 60 -190 1140
rect 3120 60 3190 1140
rect 6500 60 6570 1140
rect 9880 60 9950 1140
rect -290 -7380 -190 -6300
rect 3120 -7380 3190 -6300
rect 6500 -7380 6570 -6300
rect 9880 -7380 9950 -6300
<< nsubdiffcont >>
rect 1430 60 1500 1140
rect 4810 60 4880 1140
rect 8190 60 8260 1140
rect 11570 60 11640 1140
rect 1430 -7380 1500 -6300
rect 4810 -7380 4880 -6300
rect 8190 -7380 8260 -6300
rect 11570 -7380 11640 -6300
<< poly >>
rect 0 1230 1240 1480
rect 0 1200 400 1230
rect 840 1200 1240 1230
rect 1690 1230 2930 1480
rect 1690 1200 2090 1230
rect 2530 1200 2930 1230
rect 3380 1230 4620 1480
rect 3380 1200 3780 1230
rect 4220 1200 4620 1230
rect 5070 1230 6310 1480
rect 5070 1200 5470 1230
rect 5910 1200 6310 1230
rect 6760 1230 8000 1480
rect 6760 1200 7160 1230
rect 7600 1200 8000 1230
rect 8450 1230 9690 1480
rect 8450 1200 8850 1230
rect 9290 1200 9690 1230
rect 10140 1230 11380 1480
rect 10140 1200 10540 1230
rect 10980 1200 11380 1230
rect 0 -280 400 0
rect 840 -30 1240 0
rect 840 -160 1240 -140
rect 840 -230 870 -160
rect 1210 -230 1240 -160
rect 840 -280 1240 -230
rect 1690 -280 2090 0
rect 2530 -30 2930 0
rect 2530 -160 2930 -140
rect 2530 -230 2560 -160
rect 2900 -230 2930 -160
rect 2530 -280 2930 -230
rect 3380 -280 3780 0
rect 4220 -30 4620 0
rect 4220 -160 4620 -140
rect 4220 -230 4250 -160
rect 4590 -230 4620 -160
rect 4220 -280 4620 -230
rect 5070 -280 5470 0
rect 5910 -30 6310 0
rect 5910 -160 6310 -140
rect 5910 -230 5940 -160
rect 6280 -230 6310 -160
rect 5910 -280 6310 -230
rect 6760 -280 7160 0
rect 7600 -30 8000 0
rect 7600 -160 8000 -140
rect 7600 -230 7630 -160
rect 7970 -230 8000 -160
rect 7600 -280 8000 -230
rect 8450 -280 8850 0
rect 9290 -30 9690 0
rect 9290 -160 9690 -140
rect 9290 -230 9320 -160
rect 9660 -230 9690 -160
rect 9290 -280 9690 -230
rect 10140 -280 10540 0
rect 10980 -30 11380 0
rect 10980 -160 11380 -140
rect 10980 -230 11010 -160
rect 11350 -230 11380 -160
rect 10980 -280 11380 -230
rect 0 -1510 400 -1480
rect 840 -1510 1240 -1480
rect 1690 -1510 2090 -1480
rect 2530 -1510 2930 -1480
rect 3380 -1510 3780 -1480
rect 4220 -1510 4620 -1480
rect 5070 -1510 5470 -1480
rect 5910 -1510 6310 -1480
rect 6760 -1510 7160 -1480
rect 7600 -1510 8000 -1480
rect 8450 -1510 8850 -1480
rect 9290 -1510 9690 -1480
rect 10140 -1510 10540 -1480
rect 10980 -1510 11380 -1480
rect -630 -1830 11820 -1720
rect 0 -1860 400 -1830
rect 840 -1860 1240 -1830
rect 1690 -1860 2090 -1830
rect 2530 -1860 2930 -1830
rect 3380 -1860 3780 -1830
rect 4220 -1860 4620 -1830
rect 5070 -1860 5470 -1830
rect 5910 -1860 6310 -1830
rect 6760 -1860 7160 -1830
rect 7600 -1860 8000 -1830
rect 8450 -1860 8850 -1830
rect 9290 -1860 9690 -1830
rect 10140 -1860 10540 -1830
rect 10980 -1860 11380 -1830
rect 11420 -1860 11820 -1830
rect 0 -3090 400 -3060
rect 840 -3090 1240 -3060
rect 1690 -3090 2090 -3060
rect 2530 -3090 2930 -3060
rect 3380 -3090 3780 -3060
rect 4220 -3090 4620 -3060
rect 5070 -3090 5470 -3060
rect 5910 -3090 6310 -3060
rect 6760 -3090 7160 -3060
rect 7600 -3090 8000 -3060
rect 8450 -3090 8850 -3060
rect 9290 -3090 9690 -3060
rect 10140 -3090 10540 -3060
rect 10980 -3090 11380 -3060
rect 11420 -3090 11820 -3060
rect 0 -3180 400 -3150
rect 840 -3180 1240 -3150
rect 1690 -3180 2090 -3150
rect 2530 -3180 2930 -3150
rect 3380 -3180 3780 -3150
rect 4220 -3180 4620 -3150
rect 5070 -3180 5470 -3150
rect 5910 -3180 6310 -3150
rect 6760 -3180 7160 -3150
rect 7600 -3180 8000 -3150
rect 8450 -3180 8850 -3150
rect 9290 -3180 9690 -3150
rect 10140 -3180 10540 -3150
rect 10980 -3180 11380 -3150
rect 11420 -3180 11820 -3150
rect 0 -4410 400 -4380
rect 840 -4410 1240 -4380
rect 1690 -4410 2090 -4380
rect 2530 -4410 2930 -4380
rect 3380 -4410 3780 -4380
rect 4220 -4410 4620 -4380
rect 5070 -4410 5470 -4380
rect 5910 -4410 6310 -4380
rect 6760 -4410 7160 -4380
rect 7600 -4410 8000 -4380
rect 8450 -4410 8850 -4380
rect 9290 -4410 9690 -4380
rect 10140 -4410 10540 -4380
rect 10980 -4410 11380 -4380
rect 11420 -4410 11820 -4380
rect -630 -4520 11820 -4410
rect 0 -4760 400 -4730
rect 840 -4760 1240 -4730
rect 1690 -4760 2090 -4730
rect 2530 -4760 2930 -4730
rect 3380 -4760 3780 -4730
rect 4220 -4760 4620 -4730
rect 5070 -4760 5470 -4730
rect 5910 -4760 6310 -4730
rect 6760 -4760 7160 -4730
rect 7600 -4760 8000 -4730
rect 8450 -4760 8850 -4730
rect 9290 -4760 9690 -4730
rect 10140 -4760 10540 -4730
rect 10980 -4760 11380 -4730
rect 0 -6240 400 -5960
rect 840 -6010 1240 -5960
rect 840 -6080 870 -6010
rect 1210 -6080 1240 -6010
rect 840 -6100 1240 -6080
rect 840 -6240 1240 -6210
rect 1690 -6240 2090 -5960
rect 2530 -6010 2930 -5960
rect 2530 -6080 2560 -6010
rect 2900 -6080 2930 -6010
rect 2530 -6100 2930 -6080
rect 2530 -6240 2930 -6210
rect 3380 -6240 3780 -5960
rect 4220 -6010 4620 -5960
rect 4220 -6080 4250 -6010
rect 4590 -6080 4620 -6010
rect 4220 -6100 4620 -6080
rect 4220 -6240 4620 -6210
rect 5070 -6240 5470 -5960
rect 5910 -6010 6310 -5960
rect 5910 -6080 5940 -6010
rect 6280 -6080 6310 -6010
rect 5910 -6100 6310 -6080
rect 5910 -6240 6310 -6210
rect 6760 -6240 7160 -5960
rect 7600 -6010 8000 -5960
rect 7600 -6080 7630 -6010
rect 7970 -6080 8000 -6010
rect 7600 -6100 8000 -6080
rect 7600 -6240 8000 -6210
rect 8450 -6240 8850 -5960
rect 9290 -6010 9690 -5960
rect 9290 -6080 9320 -6010
rect 9660 -6080 9690 -6010
rect 9290 -6100 9690 -6080
rect 9290 -6240 9690 -6210
rect 10140 -6240 10540 -5960
rect 10980 -6010 11380 -5960
rect 10980 -6080 11010 -6010
rect 11350 -6080 11380 -6010
rect 10980 -6100 11380 -6080
rect 10980 -6240 11380 -6210
rect 0 -7470 400 -7440
rect 840 -7470 1240 -7440
rect 0 -7720 1240 -7470
rect 1690 -7470 2090 -7440
rect 2530 -7470 2930 -7440
rect 1690 -7720 2930 -7470
rect 3380 -7470 3780 -7440
rect 4220 -7470 4620 -7440
rect 3380 -7720 4620 -7470
rect 5070 -7470 5470 -7440
rect 5910 -7470 6310 -7440
rect 5070 -7720 6310 -7470
rect 6760 -7470 7160 -7440
rect 7600 -7470 8000 -7440
rect 6760 -7720 8000 -7470
rect 8450 -7470 8850 -7440
rect 9290 -7470 9690 -7440
rect 8450 -7720 9690 -7470
rect 10140 -7470 10540 -7440
rect 10980 -7470 11380 -7440
rect 10140 -7720 11380 -7470
<< polycont >>
rect 870 -230 1210 -160
rect 2560 -230 2900 -160
rect 4250 -230 4590 -160
rect 5940 -230 6280 -160
rect 7630 -230 7970 -160
rect 9320 -230 9660 -160
rect 11010 -230 11350 -160
rect 870 -6080 1210 -6010
rect 2560 -6080 2900 -6010
rect 4250 -6080 4590 -6010
rect 5940 -6080 6280 -6010
rect 7630 -6080 7970 -6010
rect 9320 -6080 9660 -6010
rect 11010 -6080 11350 -6010
<< locali >>
rect -310 1140 -30 1170
rect -310 60 -290 1140
rect -190 60 -130 1140
rect -60 60 -30 1140
rect -310 30 -30 60
rect 430 1130 810 1160
rect 430 60 460 1130
rect 530 60 710 1130
rect 780 60 810 1130
rect 430 -50 810 60
rect 1270 1140 1660 1170
rect 1270 60 1300 1140
rect 1370 60 1430 1140
rect 1500 60 1560 1140
rect 1630 60 1660 1140
rect 1270 30 1660 60
rect 2120 1130 2500 1160
rect 2120 60 2150 1130
rect 2220 60 2400 1130
rect 2470 60 2500 1130
rect 2120 -50 2500 60
rect 2960 1140 3350 1170
rect 2960 60 2990 1140
rect 3060 60 3120 1140
rect 3190 60 3250 1140
rect 3320 60 3350 1140
rect 2960 30 3350 60
rect 3810 1130 4190 1160
rect 3810 60 3840 1130
rect 3910 60 4090 1130
rect 4160 60 4190 1130
rect 3810 -50 4190 60
rect 4650 1140 5040 1170
rect 4650 60 4680 1140
rect 4750 60 4810 1140
rect 4880 60 4940 1140
rect 5010 60 5040 1140
rect 4650 30 5040 60
rect 5500 1130 5880 1160
rect 5500 60 5530 1130
rect 5600 60 5780 1130
rect 5850 60 5880 1130
rect 5500 -50 5880 60
rect 6340 1140 6730 1170
rect 6340 60 6370 1140
rect 6440 60 6500 1140
rect 6570 60 6630 1140
rect 6700 60 6730 1140
rect 6340 30 6730 60
rect 7190 1130 7570 1160
rect 7190 60 7220 1130
rect 7290 60 7470 1130
rect 7540 60 7570 1130
rect 7190 -50 7570 60
rect 8030 1140 8420 1170
rect 8030 60 8060 1140
rect 8130 60 8190 1140
rect 8260 60 8320 1140
rect 8390 60 8420 1140
rect 8030 30 8420 60
rect 8880 1130 9260 1160
rect 8880 60 8910 1130
rect 8980 60 9160 1130
rect 9230 60 9260 1130
rect 8880 -50 9260 60
rect 9720 1140 10110 1170
rect 9720 60 9750 1140
rect 9820 60 9880 1140
rect 9950 60 10010 1140
rect 10080 60 10110 1140
rect 9720 30 10110 60
rect 10570 1130 10950 1160
rect 10570 60 10600 1130
rect 10670 60 10850 1130
rect 10920 60 10950 1130
rect 10570 -50 10950 60
rect 11410 1140 11670 1170
rect 11410 60 11440 1140
rect 11510 60 11570 1140
rect 11640 60 11670 1140
rect 11410 30 11670 60
rect 430 -160 1240 -50
rect 430 -230 870 -160
rect 1210 -230 1240 -160
rect 430 -250 1240 -230
rect 2120 -160 2930 -50
rect 2120 -230 2560 -160
rect 2900 -230 2930 -160
rect 2120 -250 2930 -230
rect 3810 -160 4620 -50
rect 3810 -230 4250 -160
rect 4590 -230 4620 -160
rect 3810 -250 4620 -230
rect 5500 -160 6310 -50
rect 5500 -230 5940 -160
rect 6280 -230 6310 -160
rect 5500 -250 6310 -230
rect 7190 -160 8000 -50
rect 7190 -230 7630 -160
rect 7970 -230 8000 -160
rect 7190 -250 8000 -230
rect 8880 -160 9690 -50
rect 8880 -230 9320 -160
rect 9660 -230 9690 -160
rect 8880 -250 9690 -230
rect 10570 -160 11380 -50
rect 10570 -230 11010 -160
rect 11350 -230 11380 -160
rect 10570 -250 11380 -230
rect -140 -320 -20 -300
rect -140 -1440 -120 -320
rect -40 -1440 -20 -320
rect -140 -1460 -20 -1440
rect 430 -340 810 -310
rect 430 -1420 460 -340
rect 780 -1420 810 -340
rect 430 -1520 810 -1420
rect 1260 -320 1380 -300
rect 1260 -1440 1280 -320
rect 1360 -1440 1380 -320
rect 1260 -1460 1380 -1440
rect 1550 -320 1670 -300
rect 1550 -1440 1570 -320
rect 1650 -1440 1670 -320
rect 1550 -1460 1670 -1440
rect 2120 -340 2500 -310
rect 2120 -1420 2150 -340
rect 2470 -1420 2500 -340
rect 2120 -1520 2500 -1420
rect 2950 -320 3070 -300
rect 2950 -1440 2970 -320
rect 3050 -1440 3070 -320
rect 2950 -1460 3070 -1440
rect 3240 -320 3360 -300
rect 3240 -1440 3260 -320
rect 3340 -1440 3360 -320
rect 3240 -1460 3360 -1440
rect 3810 -340 4190 -310
rect 3810 -1420 3840 -340
rect 4160 -1420 4190 -340
rect 3810 -1520 4190 -1420
rect 4640 -320 4760 -300
rect 4640 -1440 4660 -320
rect 4740 -1440 4760 -320
rect 4640 -1460 4760 -1440
rect 4930 -320 5050 -300
rect 4930 -1440 4950 -320
rect 5030 -1440 5050 -320
rect 4930 -1460 5050 -1440
rect 5500 -340 5880 -310
rect 5500 -1420 5530 -340
rect 5850 -1420 5880 -340
rect 5500 -1520 5880 -1420
rect 6330 -320 6450 -300
rect 6330 -1440 6350 -320
rect 6430 -1440 6450 -320
rect 6330 -1460 6450 -1440
rect 6620 -320 6740 -300
rect 6620 -1440 6640 -320
rect 6720 -1440 6740 -320
rect 6620 -1460 6740 -1440
rect 7190 -340 7570 -310
rect 7190 -1420 7220 -340
rect 7540 -1420 7570 -340
rect 7190 -1520 7570 -1420
rect 8020 -320 8140 -300
rect 8020 -1440 8040 -320
rect 8120 -1440 8140 -320
rect 8020 -1460 8140 -1440
rect 8310 -320 8430 -300
rect 8310 -1440 8330 -320
rect 8410 -1440 8430 -320
rect 8310 -1460 8430 -1440
rect 8880 -340 9260 -310
rect 8880 -1420 8910 -340
rect 9230 -1420 9260 -340
rect 8880 -1520 9260 -1420
rect 9710 -320 9830 -300
rect 9710 -1440 9730 -320
rect 9810 -1440 9830 -320
rect 9710 -1460 9830 -1440
rect 10000 -320 10120 -300
rect 10000 -1440 10020 -320
rect 10100 -1440 10120 -320
rect 10000 -1460 10120 -1440
rect 10570 -340 10950 -310
rect 10570 -1420 10600 -340
rect 10920 -1420 10950 -340
rect 10570 -1520 10950 -1420
rect 11400 -320 11520 -300
rect 11400 -1440 11420 -320
rect 11500 -1440 11520 -320
rect 11400 -1460 11520 -1440
rect -140 -1820 810 -1520
rect 1550 -1820 2500 -1520
rect 3240 -1820 4190 -1520
rect 4930 -1820 5880 -1520
rect 6620 -1820 7570 -1520
rect 8310 -1820 9260 -1520
rect 10000 -1820 10950 -1520
rect -140 -1900 -20 -1820
rect -140 -3020 -120 -1900
rect -40 -3020 -20 -1900
rect -140 -3040 -20 -3020
rect 430 -1910 810 -1880
rect 430 -3010 460 -1910
rect 780 -3010 810 -1910
rect 430 -3040 810 -3010
rect 1260 -1900 1380 -1880
rect 1260 -3020 1280 -1900
rect 1360 -3020 1380 -1900
rect 1260 -3040 1380 -3020
rect 1550 -1900 1670 -1820
rect 1550 -3020 1570 -1900
rect 1650 -3020 1670 -1900
rect 1550 -3040 1670 -3020
rect 2120 -1910 2500 -1880
rect 2120 -3010 2150 -1910
rect 2470 -3010 2500 -1910
rect 2120 -3040 2500 -3010
rect 2950 -1900 3070 -1880
rect 2950 -3020 2970 -1900
rect 3050 -3020 3070 -1900
rect 2950 -3040 3070 -3020
rect 3240 -1900 3360 -1820
rect 3240 -3020 3260 -1900
rect 3340 -3020 3360 -1900
rect 3240 -3040 3360 -3020
rect 3810 -1910 4190 -1880
rect 3810 -3010 3840 -1910
rect 4160 -3010 4190 -1910
rect 3810 -3040 4190 -3010
rect 4640 -1900 4760 -1880
rect 4640 -3020 4660 -1900
rect 4740 -3020 4760 -1900
rect 4640 -3040 4760 -3020
rect 4930 -1900 5050 -1820
rect 4930 -3020 4950 -1900
rect 5030 -3020 5050 -1900
rect 4930 -3040 5050 -3020
rect 5500 -1910 5880 -1880
rect 5500 -3010 5530 -1910
rect 5850 -3010 5880 -1910
rect 5500 -3040 5880 -3010
rect 6330 -1900 6450 -1880
rect 6330 -3020 6350 -1900
rect 6430 -3020 6450 -1900
rect 6330 -3040 6450 -3020
rect 6620 -1900 6740 -1820
rect 6620 -3020 6640 -1900
rect 6720 -3020 6740 -1900
rect 6620 -3040 6740 -3020
rect 7190 -1910 7570 -1880
rect 7190 -3010 7220 -1910
rect 7540 -3010 7570 -1910
rect 7190 -3040 7570 -3010
rect 8020 -1900 8140 -1880
rect 8020 -3020 8040 -1900
rect 8120 -3020 8140 -1900
rect 8020 -3040 8140 -3020
rect 8310 -1900 8430 -1820
rect 8310 -3020 8330 -1900
rect 8410 -3020 8430 -1900
rect 8310 -3040 8430 -3020
rect 8880 -1910 9260 -1880
rect 8880 -3010 8910 -1910
rect 9230 -3010 9260 -1910
rect 8880 -3040 9260 -3010
rect 9710 -1900 9830 -1880
rect 9710 -3020 9730 -1900
rect 9810 -3020 9830 -1900
rect 9710 -3040 9830 -3020
rect 10000 -1900 10120 -1820
rect 10000 -3020 10020 -1900
rect 10100 -3020 10120 -1900
rect 10000 -3040 10120 -3020
rect 10570 -1910 10950 -1880
rect 10570 -3010 10600 -1910
rect 10920 -3010 10950 -1910
rect 10570 -3040 10950 -3010
rect 11840 -1900 11960 -1880
rect 11840 -3020 11860 -1900
rect 11940 -3020 11960 -1900
rect 11840 -3040 11960 -3020
rect -140 -3220 -20 -3200
rect -140 -4340 -120 -3220
rect -40 -4340 -20 -3220
rect -140 -4420 -20 -4340
rect 430 -3230 810 -3200
rect 430 -4330 460 -3230
rect 780 -4330 810 -3230
rect 430 -4360 810 -4330
rect 1260 -3220 1380 -3200
rect 1260 -4340 1280 -3220
rect 1360 -4340 1380 -3220
rect 1260 -4360 1380 -4340
rect 1550 -3220 1670 -3200
rect 1550 -4340 1570 -3220
rect 1650 -4340 1670 -3220
rect 1550 -4420 1670 -4340
rect 2120 -3230 2500 -3200
rect 2120 -4330 2150 -3230
rect 2470 -4330 2500 -3230
rect 2120 -4360 2500 -4330
rect 2950 -3220 3070 -3200
rect 2950 -4340 2970 -3220
rect 3050 -4340 3070 -3220
rect 2950 -4360 3070 -4340
rect 3240 -3220 3360 -3200
rect 3240 -4340 3260 -3220
rect 3340 -4340 3360 -3220
rect 3240 -4420 3360 -4340
rect 3810 -3230 4190 -3200
rect 3810 -4330 3840 -3230
rect 4160 -4330 4190 -3230
rect 3810 -4360 4190 -4330
rect 4640 -3220 4760 -3200
rect 4640 -4340 4660 -3220
rect 4740 -4340 4760 -3220
rect 4640 -4360 4760 -4340
rect 4930 -3220 5050 -3200
rect 4930 -4340 4950 -3220
rect 5030 -4340 5050 -3220
rect 4930 -4420 5050 -4340
rect 5500 -3230 5880 -3200
rect 5500 -4330 5530 -3230
rect 5850 -4330 5880 -3230
rect 5500 -4360 5880 -4330
rect 6330 -3220 6450 -3200
rect 6330 -4340 6350 -3220
rect 6430 -4340 6450 -3220
rect 6330 -4360 6450 -4340
rect 6620 -3220 6740 -3200
rect 6620 -4340 6640 -3220
rect 6720 -4340 6740 -3220
rect 6620 -4420 6740 -4340
rect 7190 -3230 7570 -3200
rect 7190 -4330 7220 -3230
rect 7540 -4330 7570 -3230
rect 7190 -4360 7570 -4330
rect 8020 -3220 8140 -3200
rect 8020 -4340 8040 -3220
rect 8120 -4340 8140 -3220
rect 8020 -4360 8140 -4340
rect 8310 -3220 8430 -3200
rect 8310 -4340 8330 -3220
rect 8410 -4340 8430 -3220
rect 8310 -4420 8430 -4340
rect 8880 -3230 9260 -3200
rect 8880 -4330 8910 -3230
rect 9230 -4330 9260 -3230
rect 8880 -4360 9260 -4330
rect 9710 -3220 9830 -3200
rect 9710 -4340 9730 -3220
rect 9810 -4340 9830 -3220
rect 9710 -4360 9830 -4340
rect 10000 -3220 10120 -3200
rect 10000 -4340 10020 -3220
rect 10100 -4340 10120 -3220
rect 10000 -4420 10120 -4340
rect 10570 -3230 10950 -3200
rect 10570 -4330 10600 -3230
rect 10920 -4330 10950 -3230
rect 10570 -4360 10950 -4330
rect 11840 -3220 11960 -3200
rect 11840 -4340 11860 -3220
rect 11940 -4340 11960 -3220
rect 11840 -4360 11960 -4340
rect -140 -4720 810 -4420
rect 1550 -4720 2500 -4420
rect 3240 -4720 4190 -4420
rect 4930 -4720 5880 -4420
rect 6620 -4720 7570 -4420
rect 8310 -4720 9260 -4420
rect 10000 -4720 10950 -4420
rect -140 -4800 -20 -4780
rect -140 -5920 -120 -4800
rect -40 -5920 -20 -4800
rect -140 -5940 -20 -5920
rect 430 -4820 810 -4720
rect 430 -5900 460 -4820
rect 780 -5900 810 -4820
rect 430 -5930 810 -5900
rect 1260 -4800 1380 -4780
rect 1260 -5920 1280 -4800
rect 1360 -5920 1380 -4800
rect 1260 -5940 1380 -5920
rect 1550 -4800 1670 -4780
rect 1550 -5920 1570 -4800
rect 1650 -5920 1670 -4800
rect 1550 -5940 1670 -5920
rect 2120 -4820 2500 -4720
rect 2120 -5900 2150 -4820
rect 2470 -5900 2500 -4820
rect 2120 -5930 2500 -5900
rect 2950 -4800 3070 -4780
rect 2950 -5920 2970 -4800
rect 3050 -5920 3070 -4800
rect 2950 -5940 3070 -5920
rect 3240 -4800 3360 -4780
rect 3240 -5920 3260 -4800
rect 3340 -5920 3360 -4800
rect 3240 -5940 3360 -5920
rect 3810 -4820 4190 -4720
rect 3810 -5900 3840 -4820
rect 4160 -5900 4190 -4820
rect 3810 -5930 4190 -5900
rect 4640 -4800 4760 -4780
rect 4640 -5920 4660 -4800
rect 4740 -5920 4760 -4800
rect 4640 -5940 4760 -5920
rect 4930 -4800 5050 -4780
rect 4930 -5920 4950 -4800
rect 5030 -5920 5050 -4800
rect 4930 -5940 5050 -5920
rect 5500 -4820 5880 -4720
rect 5500 -5900 5530 -4820
rect 5850 -5900 5880 -4820
rect 5500 -5930 5880 -5900
rect 6330 -4800 6450 -4780
rect 6330 -5920 6350 -4800
rect 6430 -5920 6450 -4800
rect 6330 -5940 6450 -5920
rect 6620 -4800 6740 -4780
rect 6620 -5920 6640 -4800
rect 6720 -5920 6740 -4800
rect 6620 -5940 6740 -5920
rect 7190 -4820 7570 -4720
rect 7190 -5900 7220 -4820
rect 7540 -5900 7570 -4820
rect 7190 -5930 7570 -5900
rect 8020 -4800 8140 -4780
rect 8020 -5920 8040 -4800
rect 8120 -5920 8140 -4800
rect 8020 -5940 8140 -5920
rect 8310 -4800 8430 -4780
rect 8310 -5920 8330 -4800
rect 8410 -5920 8430 -4800
rect 8310 -5940 8430 -5920
rect 8880 -4820 9260 -4720
rect 8880 -5900 8910 -4820
rect 9230 -5900 9260 -4820
rect 8880 -5930 9260 -5900
rect 9710 -4800 9830 -4780
rect 9710 -5920 9730 -4800
rect 9810 -5920 9830 -4800
rect 9710 -5940 9830 -5920
rect 10000 -4800 10120 -4780
rect 10000 -5920 10020 -4800
rect 10100 -5920 10120 -4800
rect 10000 -5940 10120 -5920
rect 10570 -4820 10950 -4720
rect 10570 -5900 10600 -4820
rect 10920 -5900 10950 -4820
rect 10570 -5930 10950 -5900
rect 11400 -4800 11520 -4780
rect 11400 -5920 11420 -4800
rect 11500 -5920 11520 -4800
rect 11400 -5940 11520 -5920
rect 430 -6010 1240 -5990
rect 430 -6080 870 -6010
rect 1210 -6080 1240 -6010
rect 430 -6190 1240 -6080
rect 2120 -6010 2930 -5990
rect 2120 -6080 2560 -6010
rect 2900 -6080 2930 -6010
rect 2120 -6190 2930 -6080
rect 3810 -6010 4620 -5990
rect 3810 -6080 4250 -6010
rect 4590 -6080 4620 -6010
rect 3810 -6190 4620 -6080
rect 5500 -6010 6310 -5990
rect 5500 -6080 5940 -6010
rect 6280 -6080 6310 -6010
rect 5500 -6190 6310 -6080
rect 7190 -6010 8000 -5990
rect 7190 -6080 7630 -6010
rect 7970 -6080 8000 -6010
rect 7190 -6190 8000 -6080
rect 8880 -6010 9690 -5990
rect 8880 -6080 9320 -6010
rect 9660 -6080 9690 -6010
rect 8880 -6190 9690 -6080
rect 10570 -6010 11380 -5990
rect 10570 -6080 11010 -6010
rect 11350 -6080 11380 -6010
rect 10570 -6190 11380 -6080
rect -310 -6300 -30 -6270
rect -310 -7380 -290 -6300
rect -190 -7380 -130 -6300
rect -60 -7380 -30 -6300
rect -310 -7410 -30 -7380
rect 430 -6300 810 -6190
rect 430 -7370 460 -6300
rect 530 -7370 710 -6300
rect 780 -7370 810 -6300
rect 430 -7400 810 -7370
rect 1270 -6300 1660 -6270
rect 1270 -7380 1300 -6300
rect 1370 -7380 1430 -6300
rect 1500 -7380 1560 -6300
rect 1630 -7380 1660 -6300
rect 1270 -7410 1660 -7380
rect 2120 -6300 2500 -6190
rect 2120 -7370 2150 -6300
rect 2220 -7370 2400 -6300
rect 2470 -7370 2500 -6300
rect 2120 -7400 2500 -7370
rect 2960 -6300 3350 -6270
rect 2960 -7380 2990 -6300
rect 3060 -7380 3120 -6300
rect 3190 -7380 3250 -6300
rect 3320 -7380 3350 -6300
rect 2960 -7410 3350 -7380
rect 3810 -6300 4190 -6190
rect 3810 -7370 3840 -6300
rect 3910 -7370 4090 -6300
rect 4160 -7370 4190 -6300
rect 3810 -7400 4190 -7370
rect 4650 -6300 5040 -6270
rect 4650 -7380 4680 -6300
rect 4750 -7380 4810 -6300
rect 4880 -7380 4940 -6300
rect 5010 -7380 5040 -6300
rect 4650 -7410 5040 -7380
rect 5500 -6300 5880 -6190
rect 5500 -7370 5530 -6300
rect 5600 -7370 5780 -6300
rect 5850 -7370 5880 -6300
rect 5500 -7400 5880 -7370
rect 6340 -6300 6730 -6270
rect 6340 -7380 6370 -6300
rect 6440 -7380 6500 -6300
rect 6570 -7380 6630 -6300
rect 6700 -7380 6730 -6300
rect 6340 -7410 6730 -7380
rect 7190 -6300 7570 -6190
rect 7190 -7370 7220 -6300
rect 7290 -7370 7470 -6300
rect 7540 -7370 7570 -6300
rect 7190 -7400 7570 -7370
rect 8030 -6300 8420 -6270
rect 8030 -7380 8060 -6300
rect 8130 -7380 8190 -6300
rect 8260 -7380 8320 -6300
rect 8390 -7380 8420 -6300
rect 8030 -7410 8420 -7380
rect 8880 -6300 9260 -6190
rect 8880 -7370 8910 -6300
rect 8980 -7370 9160 -6300
rect 9230 -7370 9260 -6300
rect 8880 -7400 9260 -7370
rect 9720 -6300 10110 -6270
rect 9720 -7380 9750 -6300
rect 9820 -7380 9880 -6300
rect 9950 -7380 10010 -6300
rect 10080 -7380 10110 -6300
rect 9720 -7410 10110 -7380
rect 10570 -6300 10950 -6190
rect 10570 -7370 10600 -6300
rect 10670 -7370 10850 -6300
rect 10920 -7370 10950 -6300
rect 10570 -7400 10950 -7370
rect 11410 -6300 11670 -6270
rect 11410 -7380 11440 -6300
rect 11510 -7380 11570 -6300
rect 11640 -7380 11670 -6300
rect 11410 -7410 11670 -7380
<< viali >>
rect -290 60 -190 1140
rect 1430 60 1500 1140
rect 3120 60 3190 1140
rect 4810 60 4880 1140
rect 6500 60 6570 1140
rect 8190 60 8260 1140
rect 9880 60 9950 1140
rect 11570 60 11640 1140
rect -120 -1440 -40 -320
rect 1280 -1440 1360 -320
rect 1570 -1440 1650 -320
rect 2970 -1440 3050 -320
rect 3260 -1440 3340 -320
rect 4660 -1440 4740 -320
rect 4950 -1440 5030 -320
rect 6350 -1440 6430 -320
rect 6640 -1440 6720 -320
rect 8040 -1440 8120 -320
rect 8330 -1440 8410 -320
rect 9730 -1440 9810 -320
rect 10020 -1440 10100 -320
rect 11420 -1440 11500 -320
rect 460 -3010 780 -1910
rect 1280 -3020 1360 -1900
rect 2150 -3010 2470 -1910
rect 2970 -3020 3050 -1900
rect 3840 -3010 4160 -1910
rect 4660 -3020 4740 -1900
rect 5530 -3010 5850 -1910
rect 6350 -3020 6430 -1900
rect 7220 -3010 7540 -1910
rect 8040 -3020 8120 -1900
rect 8910 -3010 9230 -1910
rect 9730 -3020 9810 -1900
rect 10600 -3010 10920 -1910
rect 11860 -3020 11940 -1900
rect 460 -4330 780 -3230
rect 1280 -4340 1360 -3220
rect 2150 -4330 2470 -3230
rect 2970 -4340 3050 -3220
rect 3840 -4330 4160 -3230
rect 4660 -4340 4740 -3220
rect 5530 -4330 5850 -3230
rect 6350 -4340 6430 -3220
rect 7220 -4330 7540 -3230
rect 8040 -4340 8120 -3220
rect 8910 -4330 9230 -3230
rect 9730 -4340 9810 -3220
rect 10600 -4330 10920 -3230
rect 11860 -4340 11940 -3220
rect -120 -5920 -40 -4800
rect 1280 -5920 1360 -4800
rect 1570 -5920 1650 -4800
rect 2970 -5920 3050 -4800
rect 3260 -5920 3340 -4800
rect 4660 -5920 4740 -4800
rect 4950 -5920 5030 -4800
rect 6350 -5920 6430 -4800
rect 6640 -5920 6720 -4800
rect 8040 -5920 8120 -4800
rect 8330 -5920 8410 -4800
rect 9730 -5920 9810 -4800
rect 10020 -5920 10100 -4800
rect 11420 -5920 11500 -4800
rect -290 -7380 -190 -6300
rect 1430 -7380 1500 -6300
rect 3120 -7380 3190 -6300
rect 4810 -7380 4880 -6300
rect 6500 -7380 6570 -6300
rect 8190 -7380 8260 -6300
rect 9880 -7380 9950 -6300
rect 11570 -7380 11640 -6300
<< metal1 >>
rect -300 1140 -180 1150
rect -300 60 -290 1140
rect -190 60 -180 1140
rect -300 50 -180 60
rect 1420 1140 1510 1150
rect 1420 60 1430 1140
rect 1500 60 1510 1140
rect 1420 50 1510 60
rect 3110 1140 3200 1150
rect 3110 60 3120 1140
rect 3190 60 3200 1140
rect 3110 50 3200 60
rect 4800 1140 4890 1150
rect 4800 60 4810 1140
rect 4880 60 4890 1140
rect 4800 50 4890 60
rect 6490 1140 6580 1150
rect 6490 60 6500 1140
rect 6570 60 6580 1140
rect 6490 50 6580 60
rect 8180 1140 8270 1150
rect 8180 60 8190 1140
rect 8260 60 8270 1140
rect 8180 50 8270 60
rect 9870 1140 9960 1150
rect 9870 60 9880 1140
rect 9950 60 9960 1140
rect 9870 50 9960 60
rect 11560 1140 11650 1150
rect 11560 60 11570 1140
rect 11640 60 11650 1140
rect 11560 50 11650 60
rect -140 -260 11980 -60
rect -140 -320 60 -260
rect -140 -1440 -120 -320
rect -40 -1440 60 -320
rect -140 -1460 60 -1440
rect 1180 -320 1380 -300
rect 1180 -1440 1280 -320
rect 1360 -1440 1380 -320
rect 1180 -1500 1380 -1440
rect 1550 -320 1750 -260
rect 1550 -1440 1570 -320
rect 1650 -1440 1750 -320
rect 1550 -1460 1750 -1440
rect 2870 -320 3070 -300
rect 2870 -1440 2970 -320
rect 3050 -1440 3070 -320
rect 2870 -1500 3070 -1440
rect 3240 -320 3440 -260
rect 3240 -1440 3260 -320
rect 3340 -1440 3440 -320
rect 3240 -1460 3440 -1440
rect 4560 -320 4760 -300
rect 4560 -1440 4660 -320
rect 4740 -1440 4760 -320
rect 4560 -1500 4760 -1440
rect 4930 -320 5130 -260
rect 4930 -1440 4950 -320
rect 5030 -1440 5130 -320
rect 4930 -1460 5130 -1440
rect 6250 -320 6450 -300
rect 6250 -1440 6350 -320
rect 6430 -1440 6450 -320
rect 6250 -1500 6450 -1440
rect 6620 -320 6820 -260
rect 6620 -1440 6640 -320
rect 6720 -1440 6820 -320
rect 6620 -1460 6820 -1440
rect 7940 -320 8140 -300
rect 7940 -1440 8040 -320
rect 8120 -1440 8140 -320
rect 7940 -1500 8140 -1440
rect 8310 -320 8510 -260
rect 8310 -1440 8330 -320
rect 8410 -1440 8510 -320
rect 8310 -1460 8510 -1440
rect 9630 -320 9830 -300
rect 9630 -1440 9730 -320
rect 9810 -1440 9830 -320
rect 9630 -1500 9830 -1440
rect 10000 -320 10200 -260
rect 10000 -1440 10020 -320
rect 10100 -1440 10200 -320
rect 10000 -1460 10200 -1440
rect 11320 -320 11520 -300
rect 11320 -1440 11420 -320
rect 11500 -1440 11520 -320
rect 11320 -1500 11520 -1440
rect 1180 -1700 11980 -1500
rect -630 -1910 810 -1880
rect -630 -3010 460 -1910
rect 780 -3010 810 -1910
rect -630 -3040 810 -3010
rect 1260 -1900 2500 -1880
rect 1260 -3020 1280 -1900
rect 1360 -1910 2500 -1900
rect 1360 -3010 2150 -1910
rect 2470 -3010 2500 -1910
rect 1360 -3020 2500 -3010
rect 1260 -3040 2500 -3020
rect 2950 -1900 4190 -1880
rect 2950 -3020 2970 -1900
rect 3050 -1910 4190 -1900
rect 3050 -3010 3840 -1910
rect 4160 -3010 4190 -1910
rect 3050 -3020 4190 -3010
rect 2950 -3040 4190 -3020
rect 4640 -1900 5880 -1880
rect 4640 -3020 4660 -1900
rect 4740 -1910 5880 -1900
rect 4740 -3010 5530 -1910
rect 5850 -3010 5880 -1910
rect 4740 -3020 5880 -3010
rect 4640 -3040 5880 -3020
rect 6330 -1900 7570 -1880
rect 6330 -3020 6350 -1900
rect 6430 -1910 7570 -1900
rect 6430 -3010 7220 -1910
rect 7540 -3010 7570 -1910
rect 6430 -3020 7570 -3010
rect 6330 -3040 7570 -3020
rect 8020 -1900 9260 -1880
rect 8020 -3020 8040 -1900
rect 8120 -1910 9260 -1900
rect 8120 -3010 8910 -1910
rect 9230 -3010 9260 -1910
rect 8120 -3020 9260 -3010
rect 8020 -3040 9260 -3020
rect 9710 -1900 10950 -1880
rect 9710 -3020 9730 -1900
rect 9810 -1910 10950 -1900
rect 9810 -3010 10600 -1910
rect 10920 -3010 10950 -1910
rect 9810 -3020 10950 -3010
rect 9710 -3040 10950 -3020
rect 11760 -1900 11960 -1700
rect 11760 -3020 11860 -1900
rect 11940 -3020 11960 -1900
rect 11760 -3040 11960 -3020
rect -630 -3230 810 -3200
rect -630 -4330 460 -3230
rect 780 -4330 810 -3230
rect -630 -4360 810 -4330
rect 1260 -3220 2500 -3200
rect 1260 -4340 1280 -3220
rect 1360 -3230 2500 -3220
rect 1360 -4330 2150 -3230
rect 2470 -4330 2500 -3230
rect 1360 -4340 2500 -4330
rect 1260 -4360 2500 -4340
rect 2950 -3220 4190 -3200
rect 2950 -4340 2970 -3220
rect 3050 -3230 4190 -3220
rect 3050 -4330 3840 -3230
rect 4160 -4330 4190 -3230
rect 3050 -4340 4190 -4330
rect 2950 -4360 4190 -4340
rect 4640 -3220 5880 -3200
rect 4640 -4340 4660 -3220
rect 4740 -3230 5880 -3220
rect 4740 -4330 5530 -3230
rect 5850 -4330 5880 -3230
rect 4740 -4340 5880 -4330
rect 4640 -4360 5880 -4340
rect 6330 -3220 7570 -3200
rect 6330 -4340 6350 -3220
rect 6430 -3230 7570 -3220
rect 6430 -4330 7220 -3230
rect 7540 -4330 7570 -3230
rect 6430 -4340 7570 -4330
rect 6330 -4360 7570 -4340
rect 8020 -3220 9260 -3200
rect 8020 -4340 8040 -3220
rect 8120 -3230 9260 -3220
rect 8120 -4330 8910 -3230
rect 9230 -4330 9260 -3230
rect 8120 -4340 9260 -4330
rect 8020 -4360 9260 -4340
rect 9710 -3220 10950 -3200
rect 9710 -4340 9730 -3220
rect 9810 -3230 10950 -3220
rect 9810 -4330 10600 -3230
rect 10920 -4330 10950 -3230
rect 9810 -4340 10950 -4330
rect 9710 -4360 10950 -4340
rect 11760 -3220 11960 -3200
rect 11760 -4340 11860 -3220
rect 11940 -4340 11960 -3220
rect 11760 -4540 11960 -4340
rect 1180 -4740 11980 -4540
rect -140 -4800 60 -4780
rect -140 -5920 -120 -4800
rect -40 -5920 60 -4800
rect -140 -5980 60 -5920
rect 1180 -4800 1380 -4740
rect 1180 -5920 1280 -4800
rect 1360 -5920 1380 -4800
rect 1180 -5940 1380 -5920
rect 1550 -4800 1750 -4780
rect 1550 -5920 1570 -4800
rect 1650 -5920 1750 -4800
rect 1550 -5980 1750 -5920
rect 2870 -4800 3070 -4740
rect 2870 -5920 2970 -4800
rect 3050 -5920 3070 -4800
rect 2870 -5940 3070 -5920
rect 3240 -4800 3440 -4780
rect 3240 -5920 3260 -4800
rect 3340 -5920 3440 -4800
rect 3240 -5980 3440 -5920
rect 4560 -4800 4760 -4740
rect 4560 -5920 4660 -4800
rect 4740 -5920 4760 -4800
rect 4560 -5940 4760 -5920
rect 4930 -4800 5130 -4780
rect 4930 -5920 4950 -4800
rect 5030 -5920 5130 -4800
rect 4930 -5980 5130 -5920
rect 6250 -4800 6450 -4740
rect 6250 -5920 6350 -4800
rect 6430 -5920 6450 -4800
rect 6250 -5940 6450 -5920
rect 6620 -4800 6820 -4780
rect 6620 -5920 6640 -4800
rect 6720 -5920 6820 -4800
rect 6620 -5980 6820 -5920
rect 7940 -4800 8140 -4740
rect 7940 -5920 8040 -4800
rect 8120 -5920 8140 -4800
rect 7940 -5940 8140 -5920
rect 8310 -4800 8510 -4780
rect 8310 -5920 8330 -4800
rect 8410 -5920 8510 -4800
rect 8310 -5980 8510 -5920
rect 9630 -4800 9830 -4740
rect 9630 -5920 9730 -4800
rect 9810 -5920 9830 -4800
rect 9630 -5940 9830 -5920
rect 10000 -4800 10200 -4780
rect 10000 -5920 10020 -4800
rect 10100 -5920 10200 -4800
rect 10000 -5980 10200 -5920
rect 11320 -4800 11520 -4740
rect 11320 -5920 11420 -4800
rect 11500 -5920 11520 -4800
rect 11320 -5940 11520 -5920
rect -140 -6180 11980 -5980
rect -300 -6300 -180 -6290
rect -300 -7380 -290 -6300
rect -190 -7380 -180 -6300
rect -300 -7390 -180 -7380
rect 1420 -6300 1510 -6290
rect 1420 -7380 1430 -6300
rect 1500 -7380 1510 -6300
rect 1420 -7390 1510 -7380
rect 3110 -6300 3200 -6290
rect 3110 -7380 3120 -6300
rect 3190 -7380 3200 -6300
rect 3110 -7390 3200 -7380
rect 4800 -6300 4890 -6290
rect 4800 -7380 4810 -6300
rect 4880 -7380 4890 -6300
rect 4800 -7390 4890 -7380
rect 6490 -6300 6580 -6290
rect 6490 -7380 6500 -6300
rect 6570 -7380 6580 -6300
rect 6490 -7390 6580 -7380
rect 8180 -6300 8270 -6290
rect 8180 -7380 8190 -6300
rect 8260 -7380 8270 -6300
rect 8180 -7390 8270 -7380
rect 9870 -6300 9960 -6290
rect 9870 -7380 9880 -6300
rect 9950 -7380 9960 -6300
rect 9870 -7390 9960 -7380
rect 11560 -6300 11650 -6290
rect 11560 -7380 11570 -6300
rect 11640 -7380 11650 -6300
rect 11560 -7390 11650 -7380
<< via1 >>
rect -290 60 -190 1140
rect 1430 60 1500 1140
rect 3120 60 3190 1140
rect 4810 60 4880 1140
rect 6500 60 6570 1140
rect 8190 60 8260 1140
rect 9880 60 9950 1140
rect 11570 60 11640 1140
rect -290 -7380 -190 -6300
rect 1430 -7380 1500 -6300
rect 3120 -7380 3190 -6300
rect 4810 -7380 4880 -6300
rect 6500 -7380 6570 -6300
rect 8190 -7380 8260 -6300
rect 9880 -7380 9950 -6300
rect 11570 -7380 11640 -6300
<< metal2 >>
rect 650 1260 11980 1480
rect -630 1140 590 1200
rect -630 60 -290 1140
rect -190 60 590 1140
rect -630 -60 590 60
rect 650 1140 2280 1260
rect 650 60 1430 1140
rect 1500 60 2280 1140
rect 650 0 2280 60
rect 2340 1140 3970 1200
rect 2340 60 3120 1140
rect 3190 60 3970 1140
rect 2340 -60 3970 60
rect 4030 1140 5660 1260
rect 4030 60 4810 1140
rect 4880 60 5660 1140
rect 4030 0 5660 60
rect 5720 1140 7350 1200
rect 5720 60 6500 1140
rect 6570 60 7350 1140
rect 5720 -60 7350 60
rect 7410 1140 9040 1260
rect 7410 60 8190 1140
rect 8260 60 9040 1140
rect 7410 0 9040 60
rect 9100 1140 10730 1200
rect 9100 60 9880 1140
rect 9950 60 10730 1140
rect 9100 -60 10730 60
rect -630 -280 10730 -60
rect 10790 1140 11980 1260
rect 10790 60 11570 1140
rect 11640 60 11980 1140
rect -630 -5960 590 -280
rect -630 -6180 10730 -5960
rect -630 -6300 590 -6180
rect -630 -7380 -290 -6300
rect -190 -7380 590 -6300
rect -630 -7440 590 -7380
rect 650 -6300 2280 -6240
rect 650 -7380 1430 -6300
rect 1500 -7380 2280 -6300
rect 650 -7500 2280 -7380
rect 2340 -6300 3970 -6180
rect 2340 -7380 3120 -6300
rect 3190 -7380 3970 -6300
rect 2340 -7440 3970 -7380
rect 4030 -6300 5660 -6240
rect 4030 -7380 4810 -6300
rect 4880 -7380 5660 -6300
rect 4030 -7500 5660 -7380
rect 5720 -6300 7350 -6180
rect 5720 -7380 6500 -6300
rect 6570 -7380 7350 -6300
rect 5720 -7440 7350 -7380
rect 7410 -6300 9040 -6240
rect 7410 -7380 8190 -6300
rect 8260 -7380 9040 -6300
rect 7410 -7500 9040 -7380
rect 9100 -6300 10730 -6180
rect 9100 -7380 9880 -6300
rect 9950 -7380 10730 -6300
rect 9100 -7440 10730 -7380
rect 10790 -6300 11980 60
rect 10790 -7380 11570 -6300
rect 11640 -7380 11980 -6300
rect 10790 -7500 11980 -7380
rect 650 -7720 11980 -7500
<< labels >>
rlabel metal2 -630 -6850 -630 -6850 7 Vn
port 2 w
rlabel metal2 11980 -6840 11980 -6840 3 Vp
port 1 e
rlabel poly -630 -1780 -630 -1780 7 Vg
port 4 w
rlabel metal1 -630 -2430 -630 -2430 7 Iin
port 3 w
rlabel metal1 -630 -3770 -630 -3770 7 Iin_i
port 20 w
rlabel poly -630 -4470 -630 -4470 7 Vg_i
port 19 w
rlabel poly 620 1480 620 1480 1 B6
port 5 n
rlabel poly 2320 1480 2320 1480 1 B5
port 6 n
rlabel poly 3990 1480 3990 1480 1 B4
port 7 n
rlabel poly 5690 1480 5690 1480 1 B3
port 8 n
rlabel poly 7370 1480 7370 1480 1 B2
port 9 n
rlabel poly 9070 1480 9070 1480 1 B1
port 10 n
rlabel poly 10750 1480 10750 1480 1 B0
port 11 n
rlabel metal1 11980 -1590 11980 -1590 3 Idump
port 22 e
rlabel metal1 11980 -150 11980 -150 3 Iout
port 21 e
rlabel metal1 11980 -4640 11980 -4640 3 Idump_i
port 23 e
rlabel metal1 11980 -6080 11980 -6080 3 Iout_i
port 24 e
rlabel poly 10750 -7720 10750 -7720 5 B0_i
port 18 s
rlabel poly 9070 -7720 9070 -7720 5 B1_i
port 17 s
rlabel poly 7370 -7720 7370 -7720 5 B2_i
port 16 s
rlabel poly 5700 -7720 5700 -7720 5 B3_i
port 15 s
rlabel poly 3990 -7720 3990 -7720 5 B4_i
port 14 s
rlabel poly 2320 -7720 2320 -7720 5 B5_i
port 13 s
rlabel poly 620 -7720 620 -7720 5 B6_i
port 12 s
<< end >>
