magic
tech sky130A
magscale 1 2
timestamp 1701051468
<< error_p >>
rect 1140 81 1141 2320
rect 1140 80 1260 81
rect 1140 -2619 1141 -380
rect 1140 -2620 1260 -2619
<< nwell >>
rect -1360 -2940 3760 2640
<< pmos >>
rect -1060 0 -260 2400
rect 0 0 800 2400
rect 1600 0 2400 2400
rect 2660 0 3460 2400
rect -1060 -2700 -260 -300
rect 0 -2700 800 -300
rect 1600 -2700 2400 -300
rect 2660 -2700 3460 -300
<< pdiff >>
rect -1320 2320 -1060 2400
rect -1320 80 -1240 2320
rect -1140 80 -1060 2320
rect -1320 0 -1060 80
rect -260 0 0 2400
rect 800 2320 1060 2400
rect 1340 2320 1600 2400
rect 800 80 880 2320
rect 980 80 1060 2320
rect 1340 80 1420 2320
rect 1520 80 1600 2320
rect 800 0 1060 80
rect 1340 0 1600 80
rect 2400 0 2660 2400
rect 3460 2320 3720 2400
rect 3460 80 3540 2320
rect 3640 80 3720 2320
rect 3460 0 3720 80
rect -1320 -380 -1060 -300
rect -1320 -2620 -1240 -380
rect -1140 -2620 -1060 -380
rect -1320 -2700 -1060 -2620
rect -260 -2700 0 -300
rect 800 -380 1060 -300
rect 1340 -380 1600 -300
rect 800 -2620 880 -380
rect 980 -2620 1060 -380
rect 1340 -2620 1420 -380
rect 1520 -2620 1600 -380
rect 800 -2700 1060 -2620
rect 1340 -2700 1600 -2620
rect 2400 -2700 2660 -300
rect 3460 -380 3720 -300
rect 3460 -2620 3540 -380
rect 3640 -2620 3720 -380
rect 3460 -2700 3720 -2620
<< pdiffc >>
rect -1240 80 -1140 2320
rect 880 80 980 2320
rect 1420 80 1520 2320
rect 3540 80 3640 2320
rect -1240 -2620 -1140 -380
rect 880 -2620 980 -380
rect 1420 -2620 1520 -380
rect 3540 -2620 3640 -380
<< nsubdiff >>
rect 1060 2320 1340 2400
rect 1060 80 1140 2320
rect 1260 80 1340 2320
rect 1060 0 1340 80
rect 1060 -380 1340 -300
rect 1060 -2620 1140 -380
rect 1260 -2620 1340 -380
rect 1060 -2700 1340 -2620
<< nsubdiffcont >>
rect 1140 80 1260 2320
rect 1140 -2620 1260 -380
<< poly >>
rect 0 2600 800 2640
rect 0 2500 40 2600
rect 760 2500 800 2600
rect -1060 2400 -260 2460
rect 0 2400 800 2500
rect 1600 2600 2400 2640
rect 1600 2500 1640 2600
rect 2360 2500 2400 2600
rect 1600 2400 2400 2500
rect 2660 2400 3460 2460
rect -1060 -100 -260 0
rect 0 -60 800 0
rect 1600 -60 2400 0
rect -1060 -200 -1020 -100
rect -300 -200 -260 -100
rect -1060 -300 -260 -200
rect 2660 -100 3460 0
rect 2660 -200 2700 -100
rect 3420 -200 3460 -100
rect 0 -300 800 -240
rect 1600 -300 2400 -240
rect 2660 -300 3460 -200
rect -1060 -2760 -260 -2700
rect 0 -2800 800 -2700
rect 0 -2900 40 -2800
rect 760 -2900 800 -2800
rect 0 -2940 800 -2900
rect 1600 -2800 2400 -2700
rect 2660 -2760 3460 -2700
rect 1600 -2900 1640 -2800
rect 2360 -2900 2400 -2800
rect 1600 -2940 2400 -2900
<< polycont >>
rect 40 2500 760 2600
rect 1640 2500 2360 2600
rect -1020 -200 -300 -100
rect 2700 -200 3420 -100
rect 40 -2900 760 -2800
rect 1640 -2900 2360 -2800
<< locali >>
rect -1280 2600 2400 2640
rect -1280 2500 40 2600
rect 760 2500 1640 2600
rect 2360 2500 2400 2600
rect -1280 2460 2400 2500
rect -1280 2360 -1100 2460
rect -1380 2320 -1100 2360
rect -1380 80 -1240 2320
rect -1140 80 -1100 2320
rect -1380 40 -1100 80
rect 840 2320 1560 2360
rect 840 80 880 2320
rect 980 80 1140 2320
rect 1260 80 1420 2320
rect 1520 80 1560 2320
rect 840 40 1560 80
rect 3500 2320 3780 2360
rect 3500 80 3540 2320
rect 3640 80 3780 2320
rect 3500 40 3780 80
rect -1380 -100 3780 -60
rect -1380 -200 -1020 -100
rect -300 -200 2700 -100
rect 3420 -200 3780 -100
rect -1380 -240 3780 -200
rect -1380 -380 -1100 -340
rect -1380 -2620 -1240 -380
rect -1140 -2620 -1100 -380
rect -1380 -2660 -1100 -2620
rect 840 -380 1560 -340
rect 840 -2620 880 -380
rect 980 -2620 1140 -380
rect 1260 -2620 1420 -380
rect 1520 -2620 1560 -380
rect 840 -2660 1560 -2620
rect 3500 -380 3780 -340
rect 3500 -2620 3540 -380
rect 3640 -2620 3780 -380
rect 3500 -2660 3780 -2620
rect -1280 -2760 -1100 -2660
rect -1280 -2800 2400 -2760
rect -1280 -2900 40 -2800
rect 760 -2900 1640 -2800
rect 2360 -2900 2400 -2800
rect -1280 -2940 2400 -2900
<< viali >>
rect 1140 80 1260 2320
rect 1140 -2620 1260 -380
<< metal1 >>
rect -1100 2320 3500 2640
rect -1100 80 1140 2320
rect 1260 80 3500 2320
rect -1100 -380 3500 80
rect -1100 -2620 1140 -380
rect 1260 -2620 3500 -380
rect -1100 -2760 3500 -2620
<< labels >>
rlabel locali -1380 -140 -1380 -140 7 Vcp
port 1 w
rlabel locali -1380 -1500 -1380 -1500 7 Iin1
port 3 w
rlabel locali -1380 1180 -1380 1180 7 Iin0
port 2 w
rlabel metal1 1180 2640 1180 2640 1 VP
port 4 n
rlabel locali 3780 1180 3780 1180 3 Iout0
port 5 e
rlabel locali 3780 -1500 3780 -1500 3 Iout1
port 6 e
<< end >>
