magic
tech sky130A
timestamp 1701111590
<< nwell >>
rect 710 1905 2890 5940
<< nmos >>
rect 775 515 1175 1715
rect 1320 515 1720 1715
rect 1875 515 2275 1715
rect 2420 515 2820 1715
rect 775 -880 1175 320
rect 1320 -880 1720 320
rect 1875 -880 2275 320
rect 2420 -880 2820 320
rect 890 -2275 1290 -1075
rect 1320 -2275 1720 -1075
rect 1875 -2275 2275 -1075
rect 2305 -2275 2705 -1075
<< pmos >>
rect 890 4720 1290 5920
rect 1320 4720 1720 5920
rect 1875 4720 2275 5920
rect 2305 4720 2705 5920
rect 890 3325 1290 4525
rect 1320 3325 1720 4525
rect 1875 3325 2275 4525
rect 2305 3325 2705 4525
rect 890 1930 1290 3130
rect 1320 1930 1720 3130
rect 1875 1930 2275 3130
rect 2305 1930 2705 3130
<< ndiff >>
rect 630 1655 775 1715
rect 630 575 690 1655
rect 715 575 775 1655
rect 630 515 775 575
rect 1175 1655 1320 1715
rect 1175 575 1235 1655
rect 1260 575 1320 1655
rect 1175 515 1320 575
rect 1720 1655 1875 1715
rect 1720 575 1780 1655
rect 1815 575 1875 1655
rect 1720 515 1875 575
rect 2275 1655 2420 1715
rect 2275 575 2335 1655
rect 2360 575 2420 1655
rect 2275 515 2420 575
rect 2820 1655 2965 1715
rect 2820 575 2880 1655
rect 2905 575 2965 1655
rect 2820 515 2965 575
rect 630 260 775 320
rect 630 -820 690 260
rect 715 -820 775 260
rect 630 -880 775 -820
rect 1175 260 1320 320
rect 1175 -820 1235 260
rect 1260 -820 1320 260
rect 1175 -880 1320 -820
rect 1720 260 1875 320
rect 1720 -820 1780 260
rect 1815 -820 1875 260
rect 1720 -880 1875 -820
rect 2275 260 2420 320
rect 2275 -820 2335 260
rect 2360 -820 2420 260
rect 2275 -880 2420 -820
rect 2820 260 2965 320
rect 2820 -820 2880 260
rect 2905 -820 2965 260
rect 2820 -880 2965 -820
rect 745 -1135 890 -1075
rect 745 -2215 805 -1135
rect 830 -2215 890 -1135
rect 745 -2275 890 -2215
rect 1290 -2275 1320 -1075
rect 1720 -1135 1875 -1075
rect 1720 -2215 1780 -1135
rect 1815 -2215 1875 -1135
rect 1720 -2275 1875 -2215
rect 2275 -2275 2305 -1075
rect 2705 -1135 2850 -1075
rect 2705 -2215 2765 -1135
rect 2790 -2215 2850 -1135
rect 2705 -2275 2850 -2215
<< pdiff >>
rect 745 5860 890 5920
rect 745 4780 805 5860
rect 830 4780 890 5860
rect 745 4720 890 4780
rect 1290 4720 1320 5920
rect 1720 5860 1875 5920
rect 1720 4780 1780 5860
rect 1815 4780 1875 5860
rect 1720 4720 1875 4780
rect 2275 4720 2305 5920
rect 2705 5860 2850 5920
rect 2705 4780 2765 5860
rect 2790 4780 2850 5860
rect 2705 4720 2850 4780
rect 745 4465 890 4525
rect 745 3385 805 4465
rect 830 3385 890 4465
rect 745 3325 890 3385
rect 1290 3325 1320 4525
rect 1720 4465 1875 4525
rect 1720 3385 1780 4465
rect 1815 3385 1875 4465
rect 1720 3325 1875 3385
rect 2275 3325 2305 4525
rect 2705 4465 2850 4525
rect 2705 3385 2765 4465
rect 2790 3385 2850 4465
rect 2705 3325 2850 3385
rect 745 3070 890 3130
rect 745 1990 805 3070
rect 830 1990 890 3070
rect 745 1930 890 1990
rect 1290 1930 1320 3130
rect 1720 3070 1875 3130
rect 1720 1990 1780 3070
rect 1815 1990 1875 3070
rect 1720 1930 1875 1990
rect 2275 1930 2305 3130
rect 2705 3070 2850 3130
rect 2705 1990 2765 3070
rect 2790 1990 2850 3070
rect 2705 1930 2850 1990
<< ndiffc >>
rect 690 575 715 1655
rect 1235 575 1260 1655
rect 1780 575 1815 1655
rect 2335 575 2360 1655
rect 2880 575 2905 1655
rect 690 -820 715 260
rect 1235 -820 1260 260
rect 1780 -820 1815 260
rect 2335 -820 2360 260
rect 2880 -820 2905 260
rect 805 -2215 830 -1135
rect 1780 -2215 1815 -1135
rect 2765 -2215 2790 -1135
<< pdiffc >>
rect 805 4780 830 5860
rect 1780 4780 1815 5860
rect 2765 4780 2790 5860
rect 805 3385 830 4465
rect 1780 3385 1815 4465
rect 2765 3385 2790 4465
rect 805 1990 830 3070
rect 1780 1990 1815 3070
rect 2765 1990 2790 3070
<< psubdiff >>
rect 1745 455 1850 485
rect 1745 385 1770 455
rect 1825 385 1850 455
rect 1745 350 1850 385
rect 1745 -940 1850 -910
rect 1745 -1010 1770 -940
rect 1825 -1010 1850 -940
rect 1745 -1045 1850 -1010
<< nsubdiff >>
rect 1740 4660 1855 4690
rect 1740 4590 1770 4660
rect 1825 4590 1855 4660
rect 1740 4555 1855 4590
rect 1740 3265 1855 3295
rect 1740 3195 1770 3265
rect 1825 3195 1855 3265
rect 1740 3160 1855 3195
<< psubdiffcont >>
rect 1770 385 1825 455
rect 1770 -1010 1825 -940
<< nsubdiffcont >>
rect 1770 4590 1825 4660
rect 1770 3195 1825 3265
<< poly >>
rect 600 5990 2275 6000
rect 600 5970 610 5990
rect 630 5970 2275 5990
rect 600 5960 2275 5970
rect 890 5920 1290 5935
rect 1320 5920 1720 5960
rect 1875 5920 2275 5960
rect 2305 5920 2705 5935
rect 890 4695 1290 4720
rect 890 4555 900 4695
rect 1280 4555 1290 4695
rect 890 4525 1290 4555
rect 1320 4525 1720 4720
rect 1875 4525 2275 4720
rect 2305 4695 2705 4720
rect 2305 4555 2315 4695
rect 2695 4555 2705 4695
rect 2305 4525 2705 4555
rect 890 3130 1290 3325
rect 1320 3130 1720 3325
rect 1875 3130 2275 3325
rect 2305 3130 2705 3325
rect 890 1910 1290 1930
rect 1320 1910 1720 1930
rect 1875 1910 2275 1930
rect 2305 1910 2705 1930
rect 643 1810 683 1820
rect 643 1790 653 1810
rect 673 1790 2821 1810
rect 643 1780 683 1790
rect 775 1715 1175 1790
rect 1320 1755 1720 1765
rect 1320 1735 1330 1755
rect 1710 1735 1720 1755
rect 1320 1715 1720 1735
rect 1875 1755 2275 1765
rect 1875 1735 1885 1755
rect 2265 1735 2275 1755
rect 1875 1715 2275 1735
rect 2420 1715 2820 1790
rect 775 320 1175 515
rect 1320 455 1720 515
rect 1875 455 2275 515
rect 1320 365 1720 375
rect 1320 345 1330 365
rect 1710 345 1720 365
rect 1875 365 2275 375
rect 1320 320 1720 345
rect 1875 345 1885 365
rect 2265 345 2275 365
rect 1875 320 2275 345
rect 2420 320 2820 515
rect 775 -910 1175 -880
rect 890 -1055 1175 -910
rect 890 -1075 1290 -1055
rect 1320 -1075 1720 -880
rect 1875 -1075 2275 -880
rect 2420 -910 2820 -880
rect 2420 -1055 2705 -910
rect 2305 -1075 2705 -1055
rect 890 -2295 1290 -2275
rect 1320 -2295 1720 -2275
rect 1875 -2295 2275 -2275
rect 2305 -2295 2705 -2275
<< polycont >>
rect 610 5970 630 5990
rect 900 4555 1280 4695
rect 2315 4555 2695 4695
rect 653 1790 673 1810
rect 1330 1735 1710 1755
rect 1885 1735 2265 1755
rect 1330 345 1710 365
rect 1885 345 2265 365
<< locali >>
rect 600 5990 640 6000
rect 600 5970 610 5990
rect 630 5970 640 5990
rect 600 5960 640 5970
rect 600 5909 688 5937
rect 652 5726 688 5909
rect 766 5908 2831 5956
rect 766 5890 860 5908
rect 2736 5890 2830 5908
rect 765 5860 860 5890
rect 652 5649 690 5726
rect 654 4730 690 5649
rect 765 4780 805 5860
rect 830 4780 860 5860
rect 765 4750 860 4780
rect 1750 5860 1845 5890
rect 1750 4780 1780 5860
rect 1815 4780 1845 5860
rect 1750 4750 1845 4780
rect 2735 5860 2830 5890
rect 2735 4780 2765 5860
rect 2790 4785 2830 5860
rect 2790 4780 3003 4785
rect 2735 4751 3003 4780
rect 654 4695 2707 4730
rect 890 4555 900 4695
rect 1280 4555 1290 4695
rect 1755 4660 1840 4675
rect 1755 4590 1770 4660
rect 1825 4590 1840 4660
rect 1755 4575 1840 4590
rect 890 4545 1290 4555
rect 2305 4555 2315 4695
rect 2695 4555 2705 4695
rect 2305 4545 2705 4555
rect 765 4465 860 4495
rect 765 3385 805 4465
rect 830 3385 860 4465
rect 765 3355 860 3385
rect 1750 4465 1845 4495
rect 1750 3385 1780 4465
rect 1815 3385 1845 4465
rect 1750 3355 1845 3385
rect 2735 4465 2830 4495
rect 2735 3385 2765 4465
rect 2790 3385 2830 4465
rect 2735 3355 2830 3385
rect 2964 4184 3003 4751
rect 1755 3265 1840 3280
rect 600 3235 683 3260
rect 665 1820 683 3235
rect 1755 3195 1770 3265
rect 1825 3195 1840 3265
rect 1755 3180 1840 3195
rect 765 3070 860 3100
rect 765 1990 805 3070
rect 830 1990 860 3070
rect 765 1865 860 1990
rect 1750 3070 1845 3100
rect 1750 1990 1780 3070
rect 1815 1990 1845 3070
rect 1750 1960 1845 1990
rect 2735 3070 2830 3100
rect 2735 1990 2765 3070
rect 2790 1990 2830 3070
rect 2735 1865 2830 1990
rect 643 1810 683 1820
rect 643 1790 653 1810
rect 673 1790 683 1810
rect 643 1780 683 1790
rect 700 1795 1400 1865
rect 643 1779 669 1780
rect 700 1715 745 1795
rect 1320 1765 1400 1795
rect 2195 1795 2895 1865
rect 2195 1765 2275 1795
rect 1320 1755 1720 1765
rect 1320 1735 1330 1755
rect 1710 1735 1720 1755
rect 1320 1725 1720 1735
rect 1875 1755 2275 1765
rect 1875 1735 1885 1755
rect 2265 1735 2275 1755
rect 1875 1725 2275 1735
rect 650 1655 745 1715
rect 2850 1715 2895 1795
rect 650 575 690 1655
rect 715 575 745 1655
rect 650 545 745 575
rect 1205 1655 1290 1685
rect 1205 575 1235 1655
rect 1260 575 1290 1655
rect 1205 515 1290 575
rect 1750 1655 1845 1685
rect 1750 575 1780 1655
rect 1815 575 1845 1655
rect 1750 545 1845 575
rect 2305 1655 2390 1685
rect 2305 575 2335 1655
rect 2360 575 2390 1655
rect 2305 515 2390 575
rect 2850 1655 2945 1715
rect 2850 575 2880 1655
rect 2905 575 2945 1655
rect 2850 545 2945 575
rect 600 495 2391 515
rect 1755 455 1840 470
rect 1755 385 1770 455
rect 1825 385 1840 455
rect 650 365 1720 375
rect 1755 370 1840 385
rect 650 345 1330 365
rect 1710 345 1720 365
rect 650 335 1720 345
rect 1875 365 2945 375
rect 1875 345 1885 365
rect 2265 345 2945 365
rect 1875 335 2945 345
rect 650 260 745 335
rect 650 -820 690 260
rect 715 -820 745 260
rect 650 -850 745 -820
rect 1205 260 1290 290
rect 1205 -820 1235 260
rect 1260 -820 1290 260
rect 1205 -880 1290 -820
rect 1750 260 1845 290
rect 1750 -820 1780 260
rect 1815 -820 1845 260
rect 1750 -850 1845 -820
rect 2305 260 2390 290
rect 2305 -820 2335 260
rect 2360 -820 2390 260
rect 2305 -880 2390 -820
rect 2850 260 2945 335
rect 2850 -820 2880 260
rect 2905 -820 2945 260
rect 2850 -850 2945 -820
rect 600 -900 2391 -880
rect 1755 -940 1840 -925
rect 1755 -1010 1770 -940
rect 1825 -1010 1840 -940
rect 1755 -1025 1840 -1010
rect 2964 -1104 3002 4184
rect 765 -1135 860 -1105
rect 765 -2215 805 -1135
rect 830 -2215 860 -1135
rect 765 -2261 860 -2215
rect 1750 -1135 1845 -1105
rect 1750 -2215 1780 -1135
rect 1815 -2215 1845 -1135
rect 1750 -2245 1845 -2215
rect 2735 -1135 3002 -1104
rect 2735 -2215 2765 -1135
rect 2790 -1138 3002 -1135
rect 2790 -2204 2830 -1138
rect 2790 -2215 2831 -2204
rect 765 -2262 1560 -2261
rect 2735 -2262 2831 -2215
rect 765 -2309 2831 -2262
rect 1991 -2310 2831 -2309
<< viali >>
rect 1780 4780 1815 5860
rect 1770 4590 1825 4660
rect 805 3385 830 4465
rect 1780 3385 1815 4465
rect 2765 3385 2790 4465
rect 1770 3195 1825 3265
rect 1780 1990 1815 3070
rect 1780 575 1815 1655
rect 1770 385 1825 455
rect 690 -820 715 260
rect 1780 -820 1815 260
rect 2880 -820 2905 260
rect 1770 -1010 1825 -940
rect 1780 -2215 1815 -1135
<< metal1 >>
rect 600 5860 2995 5890
rect 600 4780 1780 5860
rect 1815 4780 2995 5860
rect 600 4750 2995 4780
rect 895 4660 2700 4750
rect 895 4590 1770 4660
rect 1825 4590 2700 4660
rect 650 4465 865 4495
rect 650 3385 805 4465
rect 830 3385 865 4465
rect 650 3355 865 3385
rect 895 4465 2700 4590
rect 895 3385 1780 4465
rect 1815 3385 2700 4465
rect 650 260 750 3355
rect 895 3265 2700 3385
rect 2730 4465 2945 4495
rect 2730 3385 2765 4465
rect 2790 3385 2945 4465
rect 2730 3355 2945 3385
rect 895 3195 1770 3265
rect 1825 3195 2700 3265
rect 895 3070 2700 3195
rect 895 1990 1780 3070
rect 1815 1990 2700 3070
rect 895 1960 2700 1990
rect 650 -820 690 260
rect 715 -820 750 260
rect 650 -850 750 -820
rect 800 1655 2795 1685
rect 800 575 1780 1655
rect 1815 575 2795 1655
rect 800 455 2795 575
rect 800 385 1770 455
rect 1825 385 2795 455
rect 800 260 2795 385
rect 800 -820 1780 260
rect 1815 -820 2795 260
rect 800 -940 2795 -820
rect 2845 260 2945 3355
rect 2845 -820 2880 260
rect 2905 -820 2945 260
rect 2845 -850 2945 -820
rect 800 -1010 1770 -940
rect 1825 -1010 2795 -940
rect 800 -1075 2795 -1010
rect 600 -1135 2995 -1075
rect 600 -2215 1780 -1135
rect 1815 -2215 2995 -1135
rect 600 -2245 2995 -2215
<< labels >>
rlabel locali 600 5980 600 5980 7 Vbp
port 3 w
rlabel metal1 600 5318 600 5318 7 VP
port 2 w
rlabel metal1 600 -1679 600 -1679 7 VN
port 5 w
rlabel locali 600 -891 600 -891 7 Idac
port 6 w
rlabel locali 600 504 600 504 7 Idump
port 7 w
rlabel locali 3002 1847 3002 1847 3 Iout
port 4 e
rlabel locali 600 3248 600 3248 7 Vcn
port 8 w
rlabel locali 600 5926 600 5926 7 Vcp
port 1 w
<< end >>
