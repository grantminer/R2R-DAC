magic
tech sky130A
magscale 1 2
timestamp 1701150645
<< error_p >>
rect 39314 -9645 39315 -8348
rect 39314 -9646 39434 -9645
rect 39314 -11970 39315 -10106
<< poly >>
rect 35896 -3938 36702 -3936
rect 35232 -3970 36702 -3938
rect 35232 -4168 36326 -3970
rect 36668 -4168 36702 -3970
rect 35232 -4204 36702 -4168
<< polycont >>
rect 36326 -4168 36668 -3970
rect 4100 -15410 4240 -15250
rect 4100 -20770 4340 -20630
<< locali >>
rect 30610 -1166 31032 -1152
rect 30610 -1356 30626 -1166
rect 31016 -1356 31032 -1166
rect 30610 -1370 31032 -1356
rect 30682 -1432 31032 -1416
rect 30682 -1468 30692 -1432
rect 30958 -1468 31032 -1432
rect 30682 -1472 31032 -1468
rect 30682 -1476 30968 -1472
rect -3820 -2930 -2900 -2830
rect -3820 -3110 -3640 -2930
rect -3080 -3110 -2900 -2930
rect -3820 -3210 -2900 -3110
rect 36288 -3970 36702 -3936
rect 36288 -4168 36326 -3970
rect 36668 -4168 36702 -3970
rect 36288 -4204 36702 -4168
rect 2750 -6640 2880 -6630
rect 2750 -6700 2770 -6640
rect 2860 -6700 2880 -6640
rect 2750 -6710 2880 -6700
rect 30882 -6732 31032 -6718
rect 2750 -6768 4722 -6760
rect 2750 -6812 3974 -6768
rect 4710 -6812 4722 -6768
rect 2750 -6820 4722 -6812
rect 30882 -6852 30896 -6732
rect 31016 -6852 31032 -6732
rect 30882 -6866 31032 -6852
rect 35832 -9686 36794 -7366
rect 36288 -9812 36794 -9786
rect 36288 -9944 36318 -9812
rect 36662 -9944 36794 -9812
rect 36288 -9966 36794 -9944
rect 3866 -12120 4628 -12092
rect 2750 -12122 4628 -12120
rect 2750 -12158 3892 -12122
rect 4598 -12158 4628 -12122
rect 2750 -12170 4628 -12158
rect 2790 -12172 2922 -12170
rect 29864 -12468 31032 -12122
rect 35832 -12386 36794 -10066
rect 29866 -14764 30414 -12468
rect 29280 -14786 30414 -14764
rect 29280 -15148 29302 -14786
rect 29806 -15148 30414 -14786
rect 29280 -15172 30414 -15148
rect 30570 -15018 31032 -15000
rect 30570 -15158 30842 -15018
rect 31018 -15158 31032 -15018
rect 4060 -15250 4280 -15210
rect 4060 -15410 4100 -15250
rect 4240 -15410 4280 -15250
rect 4060 -15430 4280 -15410
rect 30570 -15482 31032 -15158
rect 2220 -15590 4580 -15530
rect 2220 -17790 2300 -15590
rect 2660 -17790 4140 -15590
rect 4500 -17790 4580 -15590
rect 30568 -15616 31032 -15482
rect 30568 -16066 31030 -15616
rect 30566 -16098 31030 -16066
rect 30566 -16530 31028 -16098
rect 30564 -16682 31028 -16530
rect 30564 -16950 31026 -16682
rect 2220 -18230 4580 -17790
rect 30562 -17146 31026 -16950
rect 30562 -18114 31024 -17146
rect 2220 -18250 4140 -18230
rect 2220 -20450 2300 -18250
rect 2660 -20430 4140 -18250
rect 4500 -20430 4580 -18230
rect 30560 -18180 31024 -18114
rect 30560 -18560 31022 -18180
rect 2660 -20450 4580 -20430
rect 2220 -20510 4580 -20450
rect 30558 -18730 31022 -18560
rect 4060 -20630 4380 -20590
rect 4060 -20770 4100 -20630
rect 4340 -20770 4380 -20630
rect 4060 -20810 4380 -20770
rect 30558 -21304 31020 -18730
rect 30556 -21328 31020 -21304
rect 30556 -21892 31018 -21328
rect 30554 -21920 31018 -21892
rect 30554 -23242 31016 -21920
rect 30552 -23362 31016 -23242
rect 30552 -23516 31014 -23362
rect 30550 -23728 31014 -23516
rect 29280 -23764 31014 -23728
rect 29280 -24096 29318 -23764
rect 29670 -23858 31014 -23764
rect 29670 -24096 31012 -23858
rect 29280 -24130 31012 -24096
<< viali >>
rect 30626 -1356 31016 -1166
rect 30692 -1468 30958 -1432
rect -3640 -3110 -3080 -2930
rect 36326 -4168 36668 -3970
rect 2770 -6700 2860 -6640
rect 3974 -6812 4710 -6768
rect 30896 -6852 31016 -6732
rect 36318 -9944 36662 -9812
rect 3892 -12158 4598 -12122
rect 29302 -15148 29806 -14786
rect 30842 -15158 31018 -15018
rect 4100 -15410 4240 -15250
rect 2300 -17790 2660 -15590
rect 4140 -17790 4500 -15590
rect 2300 -20450 2660 -18250
rect 4140 -20430 4500 -18230
rect 4100 -20770 4340 -20630
rect 29318 -24096 29670 -23764
<< metal1 >>
rect 3788 -920 4538 -918
rect 14558 -920 23354 -918
rect 3042 -924 8056 -920
rect 12782 -922 27100 -920
rect 9614 -924 31032 -922
rect 3042 -1166 31032 -924
rect 3042 -1356 30626 -1166
rect 31016 -1356 31032 -1166
rect 3042 -1368 31032 -1356
rect 3042 -1370 18130 -1368
rect 21752 -1370 31032 -1368
rect 3042 -1372 14962 -1370
rect 25684 -1372 28456 -1370
rect 3042 -1374 13644 -1372
rect -3700 -2930 -3020 -2890
rect -3700 -3110 -3640 -2930
rect -3080 -3110 -3020 -2930
rect -3700 -3150 -3020 -3110
rect 3042 -6630 3804 -1374
rect 8296 -1376 13644 -1374
rect 30682 -1432 30968 -1416
rect 30682 -1468 30692 -1432
rect 30958 -1468 30968 -1432
rect 30682 -1828 30968 -1468
rect 4724 -1830 30968 -1828
rect 3962 -2288 30968 -1830
rect 2750 -6640 3800 -6630
rect 2750 -6700 2770 -6640
rect 2860 -6700 3800 -6640
rect 2750 -6710 3800 -6700
rect 2750 -7008 2878 -6970
rect 2750 -9326 2782 -7008
rect 2850 -9326 2878 -7008
rect 2750 -9370 2878 -9326
rect 2750 -9604 2954 -9570
rect 2750 -10602 2784 -9604
rect 2698 -10754 2784 -10602
rect 2750 -11934 2784 -10754
rect 2920 -11934 2954 -9604
rect 2750 -11970 2954 -11934
rect 3040 -15090 3800 -6710
rect 3962 -6768 4726 -2288
rect 30784 -3526 31032 -3516
rect 30784 -3780 30796 -3526
rect 31020 -3780 31032 -3526
rect 30784 -3790 31032 -3780
rect 35820 -3790 38180 -1510
rect 36288 -3970 36702 -3936
rect 36288 -4168 36326 -3970
rect 36668 -4168 36702 -3970
rect 3962 -6812 3974 -6768
rect 4710 -6812 4726 -6768
rect 3962 -6824 4726 -6812
rect 4886 -6732 31032 -6606
rect 4886 -6852 30896 -6732
rect 31016 -6852 31032 -6732
rect 4886 -7070 31032 -6852
rect 3866 -7802 5584 -7070
rect 3866 -9508 4630 -7802
rect 3866 -12122 4628 -9508
rect 36288 -9812 36702 -4168
rect 37074 -7088 38180 -3790
rect 36288 -9944 36318 -9812
rect 36662 -9944 36702 -9812
rect 36288 -9966 36702 -9944
rect 3866 -12158 3892 -12122
rect 4598 -12158 4628 -12122
rect 3866 -12170 4628 -12158
rect 29280 -12290 30550 -11886
rect 29442 -14768 29832 -14764
rect 3020 -15210 3800 -15090
rect 29280 -14786 29832 -14768
rect 29280 -15148 29302 -14786
rect 29806 -15148 29832 -14786
rect 29280 -15170 29832 -15148
rect 3020 -15250 4280 -15210
rect 3020 -15410 4100 -15250
rect 4240 -15410 4280 -15250
rect 3020 -15430 4280 -15410
rect 2220 -15590 2760 -15530
rect 2220 -17790 2300 -15590
rect 2660 -17790 2760 -15590
rect 2220 -17850 2760 -17790
rect 2220 -18250 2760 -18170
rect 2220 -20450 2300 -18250
rect 2660 -20450 2760 -18250
rect 2220 -20510 2760 -20450
rect 3020 -20590 3800 -15430
rect 29442 -15512 29832 -15170
rect 30002 -14766 30550 -12290
rect 30002 -14768 30656 -14766
rect 30002 -15018 31032 -14768
rect 30002 -15158 30842 -15018
rect 31018 -15158 31032 -15018
rect 30002 -15170 31032 -15158
rect 30002 -15172 30656 -15170
rect 3020 -20630 4380 -20590
rect 3020 -20770 4100 -20630
rect 4340 -20770 4380 -20630
rect 3020 -20810 4380 -20770
rect 29442 -20850 29834 -15512
rect 31534 -17994 34414 -17780
rect 31534 -18210 31618 -17994
rect 34320 -18210 34414 -17994
rect 31534 -18264 34414 -18210
rect 29280 -21248 29834 -20850
rect 29280 -21250 29442 -21248
rect 29280 -23764 29712 -23728
rect 29280 -24096 29318 -23764
rect 29670 -24096 29712 -23764
rect 29280 -24130 29712 -24096
<< via1 >>
rect -3640 -3110 -3080 -2930
rect 2782 -9326 2850 -7008
rect 2784 -11934 2920 -9604
rect 30796 -3780 31020 -3526
rect 2300 -17790 2660 -15590
rect 2300 -20450 2660 -18250
rect 31618 -18210 34320 -17994
<< metal2 >>
rect -3700 -2930 -2140 -2890
rect -3700 -3110 -3640 -2930
rect -3080 -3110 -2140 -2930
rect -3700 -15530 -2140 -3110
rect 29012 -3526 31032 -3516
rect 29012 -3780 30796 -3526
rect 31020 -3780 31032 -3526
rect 29012 -3790 31032 -3780
rect 2750 -7008 2878 -6970
rect 2750 -9326 2782 -7008
rect 2850 -7130 2878 -7008
rect 2850 -8810 8260 -7130
rect 29012 -8810 29280 -3790
rect 2850 -9250 6620 -8810
rect 2850 -9326 2878 -9250
rect 2750 -9370 2878 -9326
rect 2750 -9604 4060 -9570
rect 2750 -11934 2784 -9604
rect 2920 -11934 4060 -9604
rect 2750 -11970 4060 -11934
rect -3700 -15590 2760 -15530
rect -3700 -17790 2300 -15590
rect 2660 -17790 2760 -15590
rect -3700 -18250 2760 -17790
rect -3700 -20450 2300 -18250
rect 2660 -20450 2760 -18250
rect -3700 -20510 2760 -20450
rect 31534 -17994 34420 -17938
rect 31534 -18210 31618 -17994
rect 34320 -18210 34420 -17994
rect 4064 -27332 6512 -26650
rect 31534 -27326 34420 -18210
rect 27870 -27332 34430 -27326
rect 4064 -28468 34430 -27332
rect 4064 -28474 30438 -28468
use bias_gen_resistor  bias_gen_resistor_0
timestamp 1701110497
transform 1 0 -15230 0 1 -12740
box 50 710 11410 12750
use bias_generator_cascode  bias_generator_cascode_0
timestamp 1701111668
transform 1 0 -3420 0 1 -13160
box -400 890 6170 6520
use cascode_mirror  cascode_mirror_0
timestamp 1701053371
transform 1 0 38174 0 1 -9726
box -1380 -2940 3780 2640
use ladder_7bit  ladder_7bit_0
timestamp 1701113382
transform 1 0 5320 0 1 -11770
box -1260 -15440 23960 2960
use output_sink  output_sink_0
timestamp 1701111590
transform 1 0 29832 0 1 -13290
box 1200 -4620 6006 12000
<< end >>
